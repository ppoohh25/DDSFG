//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10 (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sat Jul 20 20:11:15 2024

module romcoef_module (dout, clk, oce, ce, reset, ad);

output [47:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire [23:0] prom_inst_2_dout_w;
wire [23:0] prom_inst_3_dout_w;
wire [23:0] prom_inst_4_dout_w;
wire [23:0] prom_inst_5_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h559DDC123E617B8C94938874573101C9873CE78A23B43BB82D98FA53A3EA275B;
defparam prom_inst_0.INIT_RAM_01 = 256'h5CCA2F8BDE27679FCDF10D1F28281F0DF1CC9E6727DD8A2EC95BE363D945A904;
defparam prom_inst_0.INIT_RAM_02 = 256'h9C30BC3EB7268DEA3E89CB043359768A94968E7D634013DD9E5605AA46DA63E4;
defparam prom_inst_0.INIT_RAM_03 = 256'h18D2842CCB61ED71EB5CC42378C40842729AB8CDD9DCD6C6AD8B602CEEA757FE;
defparam prom_inst_0.INIT_RAM_04 = 256'hD0B088561BD78A34D46BF97EF96CD5358CDA1E598BB4D4EBF8FCF7E9D1B18754;
defparam prom_inst_0.INIT_RAM_05 = 256'hC7CDCBBFAA8C6534FBB86C17B951E066E357C1237BCA104C80AACBE3F1F7F3E6;
defparam prom_inst_0.INIT_RAM_06 = 256'hFE2A4E687981807562451FF0B7762BD77A14A42BAA1F8AED4696DD1B507B9EB7;
defparam prom_inst_0.INIT_RAM_07 = 256'h77CA13548AB8DDF80B14140AF8DCB7895212C87519B446CE4EC43195EF4189C8;
defparam prom_inst_0.INIT_RAM_08 = 256'h36AE1D83E0347EC0F8274C697C86877F6E533003CD8D45F39935C751D149B71C;
defparam prom_inst_0.INIT_RAM_09 = 256'h3CDA6FFA7DF667CE2B80CC0E47779EBBD0DBDDD6C6AC895E29EAA352F9962AB4;
defparam prom_inst_0.INIT_RAM_0A = 256'h8B4F0ABB63029825A82394FC5BB0FD407AABD3F10713161001E8C69C682AE494;
defparam prom_inst_0.INIT_RAM_0B = 256'h2711F1C8965A16C87111A835BA35A71070C6135893C5ED0D2330342F2109E8BE;
defparam prom_inst_0.INIT_RAM_0C = 256'h132227241701E2BA894E0ABD6708A02EB32FA20C6CC4125793C5EF0F26343935;
defparam prom_inst_0.INIT_RAM_0D = 256'h5186B0D2EBFA01FEF2DDBE97662CE99D48E98111971387F153ABFA407CB0DAFB;
defparam prom_inst_0.INIT_RAM_0E = 256'hE63F8FD614497597B0C0C7C5BAA5876130F7B56915B750E066E458C3257ECE14;
defparam prom_inst_0.INIT_RAM_0F = 256'hD351C73396F04189C7FC284B65767D7C715D4019EAB16F24D0730D9D24A21783;
defparam prom_inst_0.INIT_RAM_10 = 256'h1DC15BED75F46AD63A94E52D6CA2CFF20C1D25241A06E9C4955C1BD17D20BA4B;
defparam prom_inst_0.INIT_RAM_11 = 256'hC8915006B357F2840C8B026FD22D7FC7063C698DA8B9C2C1B7A4876233FBBB70;
defparam prom_inst_0.INIT_RAM_12 = 256'hD8C5A984561FDE9542E681139C1B92FF63BE105898CEFB1F3A4C55544A381CF6;
defparam prom_inst_0.INIT_RAM_13 = 256'h50626A6A614E320EDFA8681FCC700B9D26A61C8AEE499BE4245A87ACC7D9E1E1;
defparam prom_inst_0.INIT_RAM_14 = 256'h346B98BDD8EAF3F2E9D6BA966830F0A754F89426AE2EA51276D2246CACE31034;
defparam prom_inst_0.INIT_RAM_15 = 256'h8BE53780BFF6234762747D7C7360441FF1BA7930DD811CAE37B72D9BFF5AACF5;
defparam prom_inst_0.INIT_RAM_16 = 256'h57D64CB91C77C9115086B3D7F2040C0B02EFD3AD7F4807BD6A0EA93BC443B926;
defparam prom_inst_0.INIT_RAM_17 = 256'h9D40DA6BF372E854B81263ABEA204C708A9BA3A29885694314DD9C52FFA23DCE;
defparam prom_inst_0.INIT_RAM_18 = 256'h632AE89D49EC85169D1C91FD60B90A5190C5F1142E3F46453A270AE4B57C3BF1;
defparam prom_inst_0.INIT_RAM_19 = 256'hAE987A5323E9A75B06A841D158D54AB51770C007457AA5C8E1F1F8F6EBD7B993;
defparam prom_inst_0.INIT_RAM_1A = 256'h8290969286705129F7BD7A2DD87911A026A31781E33B8AD00D416C8EA6B6BCB9;
defparam prom_inst_0.INIT_RAM_1B = 256'hE51740607784898477604017E5AA6518C162F9870C88FB64C51C6BB0EC1F496A;
defparam prom_inst_0.INIT_RAM_1C = 256'hDD337FC2FC2D557389959993846D4C21EEB26D1EC666FC890D88FA62C21866AA;
defparam prom_inst_0.INIT_RAM_1D = 256'h70E857BE1B6FBAFC34648BA8BCC8CAC3B39A784C18DA9444EB891EAA2DA7177F;
defparam prom_inst_0.INIT_RAM_1E = 256'hA33ED059D950BE237FD11B5B92C1E602151F1F1706EBC89B6526DE8D33D064EE;
defparam prom_inst_0.INIT_RAM_1F = 256'h7C3AEF9A3DD768EF6DE34FB20C5DA5E41A476A85969F9E9481654012DA9A51FE;
defparam prom_inst_0.INIT_RAM_20 = 256'h01E2B9884D09BC66079F2EB431A40F70C9185E9BCFFA1C35454B493D290BE4B5;
defparam prom_inst_0.INIT_RAM_21 = 256'h3A3D37270FEDC38F530DBE66059B28AC27990161B7054984B7E0001725292518;
defparam prom_inst_0.INIT_RAM_22 = 256'h2C516D80898A8270563206D09149F89E3BCF5ADC55C42B88DD286BA4D4FB192E;
defparam prom_inst_0.INIT_RAM_23 = 256'hDE256398C3E6FF1017160BF7DBB5864E0DC37013AE40C848BE2C90EB3E87C7FE;
defparam prom_inst_0.INIT_RAM_24 = 256'h58C02076C30843759EBED5E3E8E4D7C1A279480ECA7E28C962F177F468D4368E;
defparam prom_inst_0.INIT_RAM_25 = 256'h9F29AA2290F653A7F1336C9BC2DFF3FF01FAEAD2B0855114CE7F27C55BE86BE6;
defparam prom_inst_0.INIT_RAM_26 = 256'hBB6709A232B937AC187BD5256DACE20E324D5E67665D4A2E0ADCA5651DCB700C;
defparam prom_inst_0.INIT_RAM_27 = 256'hB48144FEAF57F68C199D188AF353A9F73C78AAD4F40C1B201D10FBDCB4844A07;
defparam prom_inst_0.INIT_RAM_28 = 256'h927E623D0FD8984FFCA13DD059DA52C02683D621629BCAF10E222E30291A01DF;
defparam prom_inst_0.INIT_RAM_29 = 256'h5A686C685A4424FBCA8F4BFFA94AE372F875E955B71060A7E51A476A84959D9C;
defparam prom_inst_0.INIT_RAM_2A = 256'h1745698598A1A29A896E4B1FE9AB6413BA57EC78FA74E44CAA004D90CBFC2544;
defparam prom_inst_0.INIT_RAM_2B = 256'hCF1D619DD0FA1A32414743372204DDAC7331E69134CE5FE665DB48AB0658A1E0;
defparam prom_inst_0.INIT_RAM_2C = 256'h8BF85DB80B5495CDFB213D515B5D56452C0ADEAA6D26D77F1DB340C33EB01978;
defparam prom_inst_0.INIT_RAM_2D = 256'h53E064DF51BA1A71BF0440749EBFD7E6EDEADECAAC85561DDB913DE17B0C9514;
defparam prom_inst_0.INIT_RAM_2E = 256'h2FDB7F19AA32B22896FA56A8F2326A98BEDAEEF9FBF3E3CAA87C480BC5761EBD;
defparam prom_inst_0.INIT_RAM_2F = 256'h29F4B66F20C765FB870B85F75FBF1563A8E316406179888E8A7E694B25F5BC7A;
defparam prom_inst_0.INIT_RAM_30 = 256'h483213EBBA803DF19C3FD868EF6EE350B30E5FA8E81E4C718DA0AAAAA2917855;
defparam prom_inst_0.INIT_RAM_31 = 256'h979F9E9582674215DE9F5706AB48DC67E962D23A98ED397DB7E9113147555A56;
defparam prom_inst_0.INIT_RAM_32 = 256'h1E44617681847E6E56350BD89C5709B253EA78FE7AEE59BA1363AAE81C496C86;
defparam prom_inst_0.INIT_RAM_33 = 256'hE62A6597C1E1F9070D0AFDE8CAA3733BF9AE5AFE982AB332A9177CD82B75B6EE;
defparam prom_inst_0.INIT_RAM_34 = 256'hF85AB3034A88BDE90C26384040372409E5B88243FBAB51EE830E910B7CE34298;
defparam prom_inst_0.INIT_RAM_35 = 256'h60DF54C22681D31D5D95C4E9061A25282111F9D7AD793DF8AA53F38A189E1A8E;
defparam prom_inst_0.INIT_RAM_36 = 256'h25C154DE5FD746AD0A5FABED275880A0B6C3C8C3B6A0815928EEAB5F0BAD47D8;
defparam prom_inst_0.INIT_RAM_37 = 256'h530BBA61FF9420A31D8EF756ADFA3F7BAED8FA122128261A06E9C3955D1CD380;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000474F4F463318F4C791;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "ASYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h4149515A626A727A828A929AA2AAB2B9C1C9D0D8E0E7EFF6FE050C141B222A31;
defparam prom_inst_1.INIT_RAM_01 = 256'h252E38414A545D666F78828B949DA6AFB7C0C9D2DBE3ECF5FD060E171F283039;
defparam prom_inst_1.INIT_RAM_02 = 256'hE4EFF9040E19232D38424C57616B757F89939DA7B1BBC5CED8E2ECF5FF08121B;
defparam prom_inst_1.INIT_RAM_03 = 256'h7F8A96A2ADB9C4D0DBE7F2FE0914202B36414C57626D78838E99A4AFB9C4CFD9;
defparam prom_inst_1.INIT_RAM_04 = 256'hF4010E1B2834414E5A6773808C99A5B2BECAD7E3EFFB07131F2B37434F5B6773;
defparam prom_inst_1.INIT_RAM_05 = 256'h4553616F7D8B99A7B4C2D0DEEBF90614212F3C4A5764727F8C99A6B3C0CDDAE7;
defparam prom_inst_1.INIT_RAM_06 = 256'h7181909FAEBDCCDBEAF9081625344351606F7D8C9AA9B7C5D4E2F0FF0D1B2937;
defparam prom_inst_1.INIT_RAM_07 = 256'h79899AAABACADAEAFB0B1B2B3A4A5A6A7A8A99A9B9C8D8E7F706162534445362;
defparam prom_inst_1.INIT_RAM_08 = 256'h5C6D7F90A1B3C4D5E6F8091A2B3C4D5E6F8091A2B2C3D4E4F506162737485869;
defparam prom_inst_1.INIT_RAM_09 = 256'h1A2C3F516476899BAEC0D2E5F7091B2D3F5163758799ABBDCFE0F2041527394A;
defparam prom_inst_1.INIT_RAM_0A = 256'hB3C7DBEE0216293D5064778A9EB1C4D8EBFE1124384B5E718496A9BCCFE2F407;
defparam prom_inst_1.INIT_RAM_0B = 256'h283D51667B90A5B9CEE3F70C2035495E72869BAFC3D7EB0014283C5064788B9F;
defparam prom_inst_1.INIT_RAM_0C = 256'h788EA4BAD0E6FB11273D53687E94A9BFD4EAFF152A3F556A7F94A9BFD4E9FE13;
defparam prom_inst_1.INIT_RAM_0D = 256'hA3BAD1E8FF162E445B7289A0B7CEE4FB12283F566C8399AFC6DCF2091F354B61;
defparam prom_inst_1.INIT_RAM_0E = 256'hA9C2DAF20B233B536B839BB3CBE3FB132B425A728AA1B9D0E8FF172E465D748C;
defparam prom_inst_1.INIT_RAM_0F = 256'h8BA5BED8F10A243D566F89A2BBD4ED061F38516A829BB4CDE5FE172F48607991;
defparam prom_inst_1.INIT_RAM_10 = 256'h49637E98B3CDE8021D37516C86A0BAD4EF09233D57718AA4BED8F20B253F5872;
defparam prom_inst_1.INIT_RAM_11 = 256'hE1FD1935506C87A3BFDAF6112C48637E9AB5D0EB06213C57728DA8C3DEF8132E;
defparam prom_inst_1.INIT_RAM_12 = 256'h55728FACC9E6021F3C587592AECBE703203C597591ADC9E6021E3A56728EAAC5;
defparam prom_inst_1.INIT_RAM_13 = 256'hA5C3E1FF1D3B597794B2D0EE0B294764829FBDDAF715324F6D8AA7C4E1FE1B38;
defparam prom_inst_1.INIT_RAM_14 = 256'hD0EF0E2D4C6B8AA9C8E70625446381A0BFDDFC1B39587695B3D1F00E2C4A6987;
defparam prom_inst_1.INIT_RAM_15 = 256'hD6F61737577798B8D8F81838587898B8D7F71737567696B5D5F41433527291B0;
defparam prom_inst_1.INIT_RAM_16 = 256'hB8D9FB1C3E5F80A2C3E4052647698AABCCEC0D2E4F7091B1D2F31334547595B6;
defparam prom_inst_1.INIT_RAM_17 = 256'h7598BADDFF22446789ACCEF0123557799BBDDF0123456789ABCCEE1031537596;
defparam prom_inst_1.INIT_RAM_18 = 256'h0E3255799DC0E4082B4F7295B9DC002346698CB0D3F6193C5F82A5C7EA0D3052;
defparam prom_inst_1.INIT_RAM_19 = 256'h82A7CCF1163A5F84A9CDF2163B5F84A8CDF1153A5E82A6CAEE12365A7EA2C6EA;
defparam prom_inst_1.INIT_RAM_1A = 256'hD2F81E446A90B6DC01274D7398BEE4092F547A9FC4EA0F345A7FA4C9EE13385D;
defparam prom_inst_1.INIT_RAM_1B = 256'hFD254C739AC1E80F365D84ABD1F81F466C93B9E0072D537AA0C7ED13396086AC;
defparam prom_inst_1.INIT_RAM_1C = 256'h042D557DA5CEF61E466E96BEE60E365E85ADD5FD244C739BC3EA11396088AFD6;
defparam prom_inst_1.INIT_RAM_1D = 256'hE7103A638DB6DF08325B84ADD6FF28517AA3CCF51E466F98C0E9123A638BB4DC;
defparam prom_inst_1.INIT_RAM_1E = 256'hA5D0FA254F7AA4CFF9234E78A2CCF6214B759FC9F31C46709AC4ED17416A94BD;
defparam prom_inst_1.INIT_RAM_1F = 256'h3F6B96C2EE1945709CC7F31E4A75A0CBF7224D78A3CEF9244F7AA5D0FA25507A;
defparam prom_inst_1.INIT_RAM_20 = 256'hB5E10E3B6895C1EE1B4774A0CDF926527EABD7032F5B88B4E00C386490BCE713;
defparam prom_inst_1.INIT_RAM_21 = 256'h06346290BEEB194775A3D0FE2C5987B4E20F3D6A97C5F21F4C79A7D4012E5B88;
defparam prom_inst_1.INIT_RAM_22 = 256'h336291C0EF1E4D7CABDA09376695C3F2214F7EACDB09386694C3F11F4D7BAAD8;
defparam prom_inst_1.INIT_RAM_23 = 256'h3B6C9CCCFC2C5C8DBDED1D4C7CACDC0C3C6B9BCBFA2A5989B8E8174676A5D403;
defparam prom_inst_1.INIT_RAM_24 = 256'h205183B4E5174879AADB0C3D6E9FD001326394C5F5265787B8E819497AAADB0B;
defparam prom_inst_1.INIT_RAM_25 = 256'hE0134578AADC0F4173A6D80A3C6EA0D20536689ACCFE306293C5F7285A8BBDEE;
defparam prom_inst_1.INIT_RAM_26 = 256'h7CB0E4174B7EB2E5194C7FB3E6194C80B3E6194C7FB2E5184B7DB0E316487BAE;
defparam prom_inst_1.INIT_RAM_27 = 256'hF4295E92C7FC30659ACE03376BA0D4083D71A5D90D4276AADE124579ADE11549;
defparam prom_inst_1.INIT_RAM_28 = 256'h487EB4EA20558BC1F62C6297CD02386DA3D80D4378ADE2174D82B7EC21568BBF;
defparam prom_inst_1.INIT_RAM_29 = 256'h78AFE61D548BC2F82F669DD30A4177AEE41B5188BEF52B6197CE043A70A6DC12;
defparam prom_inst_1.INIT_RAM_2A = 256'h84BCF42C649CD40C447CB4EC235B93CB023A71A9E0184F87BEF62D649BD20A41;
defparam prom_inst_1.INIT_RAM_2B = 256'h6BA5DE175089C3FC356EA7E019528AC3FC356DA6DF175088C1F9326AA3DB134B;
defparam prom_inst_1.INIT_RAM_2C = 256'h2F69A4DE19538DC7013C76B0EA245E98D20C457FB9F32C66A0D9134C86BFF932;
defparam prom_inst_1.INIT_RAM_2D = 256'hCF0A4681BDF8346FAAE6215C97D20D4883BEF9346FAAE5205A95D00A4580BAF5;
defparam prom_inst_1.INIT_RAM_2E = 256'h4B87C4013D7AB6F32F6BA8E4205D99D5114D89C5013D79B5F12D69A5E01C5893;
defparam prom_inst_1.INIT_RAM_2F = 256'hA3E01E5C9AD7155290CE0B4886C3013E7BB8F63370ADEA2764A1DE1B5894D10E;
defparam prom_inst_1.INIT_RAM_30 = 256'hD7165593D211508ECD0C4A89C7064483C1003E7CBAF93775B3F12F6DABE92765;
defparam prom_inst_1.INIT_RAM_31 = 256'hE72767A7E72767A7E62666A6E52564A4E32362A2E120609FDE1D5D9CDB1A5998;
defparam prom_inst_1.INIT_RAM_32 = 256'hD4155697D8195A9BDC1D5E9EDF2061A1E22263A3E42465A5E62666A6E72767A7;
defparam prom_inst_1.INIT_RAM_33 = 256'h9CDF2163A5E7296CAEF03173B5F7397BBCFE4081C3054688C90B4C8DCF105192;
defparam prom_inst_1.INIT_RAM_34 = 256'h4185C80C4F92D5185C9FE22568ABEE3173B6F93C7EC1044689CC0E5193D5185A;
defparam prom_inst_1.INIT_RAM_35 = 256'hC3074C90D5195DA2E62A6EB2F73B7FC3074B8ED2165A9EE12569ACF03477BBFE;
defparam prom_inst_1.INIT_RAM_36 = 256'h2166ACF1377CC2074D92D71C62A7EC3176BB00458ACF14599EE2276CB1F53A7E;
defparam prom_inst_1.INIT_RAM_37 = 256'h5BA2E82F75BC034990D61C63A9EF367CC2084E95DB2167ADF3387EC40A5095DB;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000DD246BB2F94086CD14;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[23:0],dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 8;
defparam prom_inst_2.RESET_MODE = "ASYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFDFDFDFDFDFDFD;
defparam prom_inst_2.INIT_RAM_01 = 256'hFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFCFCFCFCFCFCFC;
defparam prom_inst_2.INIT_RAM_02 = 256'hF9F9F9FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFBFBFB;
defparam prom_inst_2.INIT_RAM_03 = 256'hF8F8F8F8F8F8F8F8F8F8F8F8F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9;
defparam prom_inst_2.INIT_RAM_04 = 256'hF6F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F8F8F8F8F8F8F8F8F8F8;
defparam prom_inst_2.INIT_RAM_05 = 256'hF5F5F5F5F5F5F5F5F5F5F5F5F5F5F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6;
defparam prom_inst_2.INIT_RAM_06 = 256'hF3F3F3F3F3F3F3F3F3F3F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F5F5F5F5;
defparam prom_inst_2.INIT_RAM_07 = 256'hF1F1F1F1F1F1F1F1F1F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F3F3F3F3F3F3F3;
defparam prom_inst_2.INIT_RAM_08 = 256'hEFEFEFEFEFEFEFEFEFEFF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F1F1F1F1F1F1F1;
defparam prom_inst_2.INIT_RAM_09 = 256'hEDEDEDEDEDEDEDEDEDEDEDEDEDEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFEFEFEFEF;
defparam prom_inst_2.INIT_RAM_0A = 256'hEAEAEAEAEBEBEBEBEBEBEBEBEBEBEBEBEBEBECECECECECECECECECECECECECED;
defparam prom_inst_2.INIT_RAM_0B = 256'hE8E8E8E8E8E8E8E8E8E8E8E9E9E9E9E9E9E9E9E9E9E9E9EAEAEAEAEAEAEAEAEA;
defparam prom_inst_2.INIT_RAM_0C = 256'hE5E5E5E5E5E5E5E6E6E6E6E6E6E6E6E6E6E6E6E7E7E7E7E7E7E7E7E7E7E7E7E8;
defparam prom_inst_2.INIT_RAM_0D = 256'hE2E2E2E2E2E3E3E3E3E3E3E3E3E3E3E3E4E4E4E4E4E4E4E4E4E4E4E5E5E5E5E5;
defparam prom_inst_2.INIT_RAM_0E = 256'hDFDFDFDFE0E0E0E0E0E0E0E0E0E0E0E1E1E1E1E1E1E1E1E1E1E1E2E2E2E2E2E2;
defparam prom_inst_2.INIT_RAM_0F = 256'hDCDCDCDCDCDDDDDDDDDDDDDDDDDDDDDEDEDEDEDEDEDEDEDEDEDEDFDFDFDFDFDF;
defparam prom_inst_2.INIT_RAM_10 = 256'hD9D9D9D9D9D9D9DADADADADADADADADADADBDBDBDBDBDBDBDBDBDBDCDCDCDCDC;
defparam prom_inst_2.INIT_RAM_11 = 256'hD5D5D6D6D6D6D6D6D6D6D6D7D7D7D7D7D7D7D7D7D8D8D8D8D8D8D8D8D8D8D9D9;
defparam prom_inst_2.INIT_RAM_12 = 256'hD2D2D2D2D2D2D3D3D3D3D3D3D3D3D3D4D4D4D4D4D4D4D4D4D5D5D5D5D5D5D5D5;
defparam prom_inst_2.INIT_RAM_13 = 256'hCECECECECFCFCFCFCFCFCFCFD0D0D0D0D0D0D0D0D0D1D1D1D1D1D1D1D1D1D2D2;
defparam prom_inst_2.INIT_RAM_14 = 256'hCACACBCBCBCBCBCBCBCBCCCCCCCCCCCCCCCCCCCDCDCDCDCDCDCDCDCECECECECE;
defparam prom_inst_2.INIT_RAM_15 = 256'hC6C6C7C7C7C7C7C7C7C7C8C8C8C8C8C8C8C8C9C9C9C9C9C9C9C9CACACACACACA;
defparam prom_inst_2.INIT_RAM_16 = 256'hC2C2C2C3C3C3C3C3C3C3C4C4C4C4C4C4C4C4C5C5C5C5C5C5C5C5C6C6C6C6C6C6;
defparam prom_inst_2.INIT_RAM_17 = 256'hBEBEBEBEBEBFBFBFBFBFBFBFC0C0C0C0C0C0C0C1C1C1C1C1C1C1C1C2C2C2C2C2;
defparam prom_inst_2.INIT_RAM_18 = 256'hBABABABABABABABBBBBBBBBBBBBBBCBCBCBCBCBCBCBCBDBDBDBDBDBDBDBEBEBE;
defparam prom_inst_2.INIT_RAM_19 = 256'hB5B5B5B5B6B6B6B6B6B6B6B7B7B7B7B7B7B7B8B8B8B8B8B8B8B9B9B9B9B9B9B9;
defparam prom_inst_2.INIT_RAM_1A = 256'hB0B0B1B1B1B1B1B1B2B2B2B2B2B2B2B3B3B3B3B3B3B3B4B4B4B4B4B4B4B5B5B5;
defparam prom_inst_2.INIT_RAM_1B = 256'hABACACACACACACADADADADADADADAEAEAEAEAEAEAFAFAFAFAFAFAFB0B0B0B0B0;
defparam prom_inst_2.INIT_RAM_1C = 256'hA7A7A7A7A7A7A7A8A8A8A8A8A8A9A9A9A9A9A9A9AAAAAAAAAAAAABABABABABAB;
defparam prom_inst_2.INIT_RAM_1D = 256'hA1A2A2A2A2A2A2A3A3A3A3A3A3A3A4A4A4A4A4A4A5A5A5A5A5A5A6A6A6A6A6A6;
defparam prom_inst_2.INIT_RAM_1E = 256'h9C9C9C9D9D9D9D9D9D9E9E9E9E9E9E9F9F9F9F9F9FA0A0A0A0A0A0A1A1A1A1A1;
defparam prom_inst_2.INIT_RAM_1F = 256'h97979797979898989898989999999999999A9A9A9A9A9A9B9B9B9B9B9B9C9C9C;
defparam prom_inst_2.INIT_RAM_20 = 256'h9191929292929292939393939393949494949495959595959596969696969697;
defparam prom_inst_2.INIT_RAM_21 = 256'h8C8C8C8C8C8C8D8D8D8D8D8D8E8E8E8E8E8F8F8F8F8F8F909090909091919191;
defparam prom_inst_2.INIT_RAM_22 = 256'h8686868686878787878788888888888889898989898A8A8A8A8A8A8B8B8B8B8B;
defparam prom_inst_2.INIT_RAM_23 = 256'h8080808080818181818182828282828383838383838484848484858585858586;
defparam prom_inst_2.INIT_RAM_24 = 256'h7A7A7A7A7A7B7B7B7B7B7C7C7C7C7C7D7D7D7D7D7D7E7E7E7E7E7F7F7F7F7F80;
defparam prom_inst_2.INIT_RAM_25 = 256'h7374747474747575757575767676767677777777777778787878787979797979;
defparam prom_inst_2.INIT_RAM_26 = 256'h6D6D6D6E6E6E6E6E6F6F6F6F6F70707070707171717171727272727273737373;
defparam prom_inst_2.INIT_RAM_27 = 256'h6667676767676868686869696969696A6A6A6A6A6B6B6B6B6B6C6C6C6C6C6D6D;
defparam prom_inst_2.INIT_RAM_28 = 256'h6060606061616161616262626263636363636464646464656565656566666666;
defparam prom_inst_2.INIT_RAM_29 = 256'h5959595A5A5A5A5A5B5B5B5B5C5C5C5C5C5D5D5D5D5D5E5E5E5E5F5F5F5F5F60;
defparam prom_inst_2.INIT_RAM_2A = 256'h5252525353535354545454545555555556565656565757575757585858585959;
defparam prom_inst_2.INIT_RAM_2B = 256'h4B4B4B4C4C4C4C4C4D4D4D4D4E4E4E4E4E4F4F4F4F5050505050515151515252;
defparam prom_inst_2.INIT_RAM_2C = 256'h44444444454545454646464646474747474848484848494949494A4A4A4A4A4B;
defparam prom_inst_2.INIT_RAM_2D = 256'h3C3D3D3D3D3D3E3E3E3E3F3F3F3F404040404041414141424242424343434343;
defparam prom_inst_2.INIT_RAM_2E = 256'h35353536363636363737373738383838393939393A3A3A3A3A3B3B3B3B3C3C3C;
defparam prom_inst_2.INIT_RAM_2F = 256'h2D2D2E2E2E2E2F2F2F2F30303030313131313132323232333333333434343435;
defparam prom_inst_2.INIT_RAM_30 = 256'h25262626262727272728282828292929292A2A2A2A2A2B2B2B2B2C2C2C2C2D2D;
defparam prom_inst_2.INIT_RAM_31 = 256'h1D1E1E1E1E1F1F1F1F2020202021212121222222222323232324242424252525;
defparam prom_inst_2.INIT_RAM_32 = 256'h15161616161717171718181818191919191A1A1A1A1B1B1B1B1C1C1C1C1D1D1D;
defparam prom_inst_2.INIT_RAM_33 = 256'h0D0D0E0E0E0E0F0F0F0F10101010111111111212121313131314141414151515;
defparam prom_inst_2.INIT_RAM_34 = 256'h050505060606060707070708080808090909090A0A0A0B0B0B0B0C0C0C0C0D0D;
defparam prom_inst_2.INIT_RAM_35 = 256'hFCFDFDFDFDFEFEFEFEFFFFFFFF00000001010101020202020303030304040404;
defparam prom_inst_2.INIT_RAM_36 = 256'hF4F4F4F4F5F5F5F6F6F6F6F7F7F7F7F8F8F8F9F9F9F9FAFAFAFAFBFBFBFBFCFC;
defparam prom_inst_2.INIT_RAM_37 = 256'hEBEBEBECECECEDEDEDEDEEEEEEEEEFEFEFF0F0F0F0F1F1F1F1F2F2F2F3F3F3F3;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000E8E9E9E9E9EAEAEAEB;
defparam prom_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[23:0],dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 8;
defparam prom_inst_3.RESET_MODE = "ASYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h974C02B76C21D68C41F6AB6015CA7F34E99E5308BD7227DC9146FAAF6419CE83;
defparam prom_inst_3.INIT_RAM_01 = 256'hE69C5208BD7329DE944AFFB56B20D68B41F6AC6117CC8237EDA2570DC2772DE2;
defparam prom_inst_3.INIT_RAM_02 = 256'h22D88F45FCB2681FD58B41F8AE641AD0873DF3A95F15CB8137EDA3590FC57A30;
defparam prom_inst_3.INIT_RAM_03 = 256'h48FFB66D24DC934A01B86F25DC934A01B86F25DC934A00B76E24DB9148FEB56B;
defparam prom_inst_3.INIT_RAM_04 = 256'h560EC67E36EEA55D15CD843CF4AB631BD28A41F9B0681FD78E45FDB46B22DA91;
defparam prom_inst_3.INIT_RAM_05 = 256'h4A03BC742DE69E5710C88139F2AA631BD48C44FDB56D25DE964E06BE762EE69E;
defparam prom_inst_3.INIT_RAM_06 = 256'h21DB954F08C27B35EEA8611BD48E4700B9732CE59E5711CA833CF5AE6720D891;
defparam prom_inst_3.INIT_RAM_07 = 256'hDA944F0AC47F3AF4AF6924DE98530DC7823CF6B06A24DE98520CC6803AF4AE68;
defparam prom_inst_3.INIT_RAM_08 = 256'h712DE8A4601CD7934E0AC5813CF8B36E2AE5A05B16D28D4803BE7934EFA9641F;
defparam prom_inst_3.INIT_RAM_09 = 256'hE4A15E1BD895510ECB884401BD7A36F3AF6C28E4A05D19D5914D09C5813DF9B5;
defparam prom_inst_3.INIT_RAM_0A = 256'h32F0AE6C2AE8A66422E09E5C19D7955210CD8B4806C3813EFBB97633F0AD6A27;
defparam prom_inst_3.INIT_RAM_0B = 256'h5716D6955514D3925111D08F4E0DCC8B4908C7864403C2803FFDBC7A39F7B573;
defparam prom_inst_3.INIT_RAM_0C = 256'h5112D3945415D6965717D8985919D9995A1ADA9A5A1ADA9A5A19D9995918D897;
defparam prom_inst_3.INIT_RAM_0D = 256'h1FE1A36628EAAC6E30F2B47537F9BB7C3EFFC1824405C788490ACB8D4E0FD090;
defparam prom_inst_3.INIT_RAM_0E = 256'hBD814508CC905317DA9E6124E7AB6E31F4B77A3D00C386480BCE905315D89A5D;
defparam prom_inst_3.INIT_RAM_0F = 256'h2AEFB47A3F04C98E5318DDA2672CF0B57A3E03C78C5015D99D6125E9AD7135F9;
defparam prom_inst_3.INIT_RAM_10 = 256'h6229F0B77E450CD2996026EDB37A4006CD93591FE5AB7137FDC3884E14D99F64;
defparam prom_inst_3.INIT_RAM_11 = 256'h652DF6BF875018E1A9723A02CA925A22EAB27A420AD1996128F0B77E460DD49B;
defparam prom_inst_3.INIT_RAM_12 = 256'h2EF9C38E5823EDB7814B15DFA9733D07D19A642DF7C08A531CE6AF78410AD39C;
defparam prom_inst_3.INIT_RAM_13 = 256'hBD895622EEBB87531FEBB7834E1AE6B27D4914DFAB76410CD8A36E3803CE9964;
defparam prom_inst_3.INIT_RAM_14 = 256'h0EDDAB794816E4B2804E1CE9B7855220EDBB885523F0BD8A5724F1BE8A5724F0;
defparam prom_inst_3.INIT_RAM_15 = 256'h20F0C191613202D2A2724111E1B180501FEFBE8D5D2CFBCA99683705D4A37140;
defparam prom_inst_3.INIT_RAM_16 = 256'hF0C295673A0CDEB0825426F8CA9B6D3F10E2B3855627F8C99A6B3C0DDEAE7F50;
defparam prom_inst_3.INIT_RAM_17 = 256'h7B5025F9CEA2764B1FF3C79B6F4317EBBE9265390CE0B386592CFFD2A5784B1D;
defparam prom_inst_3.INIT_RAM_18 = 256'hC0976E451CF2C99F764C22F9CFA57B5127FDD2A87E5329FED3A87E5328FDD2A7;
defparam prom_inst_3.INIT_RAM_19 = 256'hBC956F4821FAD3AB845D350EE6BF976F471FF8CFA77F572F06DEB58C643B12E9;
defparam prom_inst_3.INIT_RAM_1A = 256'h6D482400DBB6926D4823FED9B48E69441EF8D3AD87613C16EFC9A37D563009E3;
defparam prom_inst_3.INIT_RAM_1B = 256'hD0AE8C6A482603E1BF9C79573411EECBA885623F1BF8D4B18D694521FED9B591;
defparam prom_inst_3.INIT_RAM_1C = 256'hE3C4A48565462606E6C6A68665452504E4C3A28261401FFEDCBB9A78573514F2;
defparam prom_inst_3.INIT_RAM_1D = 256'hA4876B4E3114F6D9BC9E816346280AECCEB09274553718FADBBD9E7F60412202;
defparam prom_inst_3.INIT_RAM_1E = 256'h11F7DCC2A88D73583E2308EDD2B79C81654A2E13F7DBBFA3876B4F3316FADDC1;
defparam prom_inst_3.INIT_RAM_1F = 256'h260FF8E0C8B199816951392109F0D8BFA78E755C432A11F8DEC5AB92785E452B;
defparam prom_inst_3.INIT_RAM_20 = 256'hE3CEBAA5907B66513C2712FCE7D1BBA6907A644E38210BF4DEC7B19A836C553E;
defparam prom_inst_3.INIT_RAM_21 = 256'h4432210FFDEBD9C7B4A2907D6A5845321F0CF9E5D2BFAB9784705C4834200CF7;
defparam prom_inst_3.INIT_RAM_22 = 256'h47382A1B0CFDEEDFCFC0B0A191817161514131211000EFDECEBDAC9B89786755;
defparam prom_inst_3.INIT_RAM_23 = 256'hEADFD3C7BBAFA3978B7E7265584C3F3225180AFDF0E2D5C7B9AB9D8F81736456;
defparam prom_inst_3.INIT_RAM_24 = 256'h2B231A1108FFF6EDE4DBD1C8BEB5ABA1978D83796E64594F44392E23180D01F6;
defparam prom_inst_3.INIT_RAM_25 = 256'h0702FCF7F1EBE6E0DAD3CDC7C0BAB3ADA69F989189827B736C645C544C443C33;
defparam prom_inst_3.INIT_RAM_26 = 256'h7C7A787673716E6B696663605C5956524F4B47433F3B37322E2A25201B16110C;
defparam prom_inst_3.INIT_RAM_27 = 256'h88898A8B8C8D8E8E8F8F9090909090908F8F8E8E8D8C8B8A898886858382807E;
defparam prom_inst_3.INIT_RAM_28 = 256'h282D31363A3E42464A4E5255595C5F6266686B6E717376787A7C7E8082838587;
defparam prom_inst_3.INIT_RAM_29 = 256'h5A626A727A828991989FA6ADB4BBC2C9CFD5DCE2E8EEF4F9FF040A0F14191E23;
defparam prom_inst_3.INIT_RAM_2A = 256'h1C28333F4A55616C76818C96A1ABB5BFC9D3DDE7F0FA030C151E273039414A52;
defparam prom_inst_3.INIT_RAM_2B = 256'h6C7B8A99A8B7C6D4E3F1FF0E1C29374552606D7B8895A2AEBBC8D4E0EDF90510;
defparam prom_inst_3.INIT_RAM_2C = 256'h47596C7F92A4B7C9DBEDFF112234455768798A9BACBCCDDDEEFE0E1E2E3D4D5C;
defparam prom_inst_3.INIT_RAM_2D = 256'hAAC1D8EE041B31475D72889EB3C8DDF2071C31465A6E8397ABBFD2E6FA0D2033;
defparam prom_inst_3.INIT_RAM_2E = 256'h95AFC9E4FE18324C657F98B2CBE4FD162F47607890A9C1D8F0081F374E657C93;
defparam prom_inst_3.INIT_RAM_2F = 256'h0322405E7C9AB8D6F3112E4B6885A2BFDBF814304D6984A0BCD7F30E29445F7A;
defparam prom_inst_3.INIT_RAM_30 = 256'hF416395B7D9FC0E20425466789A9CAEB0B2C4C6C8CACCCEC0B2B4A6988A7C6E5;
defparam prom_inst_3.INIT_RAM_31 = 256'h648BB1D7FD23496F94BADF04294E7398BCE105294D7195B9DC002346698CAFD1;
defparam prom_inst_3.INIT_RAM_32 = 256'h527DA7D2FC26507AA3CDF61F49729AC3EC143D658DB5DD052C547BA2C9F0173E;
defparam prom_inst_3.INIT_RAM_33 = 256'hBCEA194776A4D2002E5C89B7E4113E6B98C4F11D4A76A2CDF925507CA7D2FD28;
defparam prom_inst_3.INIT_RAM_34 = 256'h9ED10436699BCE00326496C7F92A5C8DBEEF1F5080B1E1114171A0D0FF2F5E8D;
defparam prom_inst_3.INIT_RAM_35 = 256'hF72E659CD30A4177ADE41A5086BBF1265C91C6FB2F6498CD0135699DD004376B;
defparam prom_inst_3.INIT_RAM_36 = 256'hC4003B77B2ED28639ED8134D87C1FB356FA8E21B548DC6FF3770A8E0185088BF;
defparam prom_inst_3.INIT_RAM_37 = 256'h034484C3034382C201407FBEFC3B79B7F53371AFEC2A67A4E11E5B97D4104C88;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000BBFD3E7FC0014283C3;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[23:0],dout[39:32]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 8;
defparam prom_inst_4.RESET_MODE = "ASYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hB4A494837363524232211101F1E0D0C0AF9F8F7F6E5E4E3D2D1D0CFCECDCCBBB;
defparam prom_inst_4.INIT_RAM_01 = 256'hBDAD9D8D7C6C5C4B3B2B1A0AFAEAD9C9B9A898887867574736261606F5E5D5C4;
defparam prom_inst_4.INIT_RAM_02 = 256'hC7B6A696857565554434241303F3E3D2C2B2A19181716050402F1F0FFFEEDECE;
defparam prom_inst_4.INIT_RAM_03 = 256'hD0BFAF9F8F7E6E5E4E3D2D1D0CFCECDCCBBBAB9A8A7A6A594939281808F7E7D7;
defparam prom_inst_4.INIT_RAM_04 = 256'hD9C9B8A898877767574636261505F5E5D4C4B4A393837362524231211101F0E0;
defparam prom_inst_4.INIT_RAM_05 = 256'hE2D2C1B1A1908070604F3F2F1E0EFEEEDDCDBDAC9C8C7C6B5B4B3B2A1A0AF9E9;
defparam prom_inst_4.INIT_RAM_06 = 256'hEBDACABAAA99897968584838271707F7E6D6C6B5A595857464544333231302F2;
defparam prom_inst_4.INIT_RAM_07 = 256'hF3E3D3C3B2A2928171615140302010FFEFDFCEBEAE9E8D7D6D5D4C3C2C1B0BFB;
defparam prom_inst_4.INIT_RAM_08 = 256'hFCECDBCBBBAB9A8A7A6A594939281808F8E7D7C7B7A696867665554534241404;
defparam prom_inst_4.INIT_RAM_09 = 256'h04F4E4D4C3B3A393827262524131211000F0E0CFBFAF9F8E7E6E5E4D3D2D1C0C;
defparam prom_inst_4.INIT_RAM_0A = 256'h0DFCECDCCCBBAB9B8B7A6A5A4A39291909F8E8D8C8B7A7978676665645352515;
defparam prom_inst_4.INIT_RAM_0B = 256'h1505F4E4D4C4B3A393837262524231211101F0E0D0C0AF9F8F7E6E5E4E3D2D1D;
defparam prom_inst_4.INIT_RAM_0C = 256'h1D0DFCECDCCCBBAB9B8B7A6A5A4A39291909F8E8D8C8B7A79787766656463525;
defparam prom_inst_4.INIT_RAM_0D = 256'h251404F4E4D3C3B3A392827262514131211000F0E0D0BFAF9F8F7E6E5E4E3D2D;
defparam prom_inst_4.INIT_RAM_0E = 256'h2C1C0CFCEBDBCBBBAA9A8A7A69594939281808F8E8D7C7B7A796867666554535;
defparam prom_inst_4.INIT_RAM_0F = 256'h34231303F3E3D2C2B2A2918171615040302010FFEFDFCFBEAE9E8E7D6D5D4D3C;
defparam prom_inst_4.INIT_RAM_10 = 256'h3B2B1A0AFAEADAC9B9A999887868584837271707F6E6D6C6B5A5958575645444;
defparam prom_inst_4.INIT_RAM_11 = 256'h4232211101F1E1D0C0B0A0907F6F5F4F3E2E1E0EFEEDDDCDBDAC9C8C7C6C5B4B;
defparam prom_inst_4.INIT_RAM_12 = 256'h4938281808F8E7D7C7B7A796867666564535251504F4E4D4C4B3A39383736252;
defparam prom_inst_4.INIT_RAM_13 = 256'h4F3F2F1F0EFEEEDECEBDAD9D8D7D6C5C4C3C2C1B0BFBEBDBCABAAA9A8A796959;
defparam prom_inst_4.INIT_RAM_14 = 256'h564535251505F4E4D4C4B4A393837363524232221201F1E1D1C1B0A09080705F;
defparam prom_inst_4.INIT_RAM_15 = 256'h5C4B3B2B1B0BFBEADACABAAA99897969594838281808F7E7D7C7B7A796867666;
defparam prom_inst_4.INIT_RAM_16 = 256'h61514131211100F0E0D0C0AF9F8F7F6F5F4E3E2E1E0EFDEDDDCDBDAD9C8C7C6C;
defparam prom_inst_4.INIT_RAM_17 = 256'h67574736261606F6E6D5C5B5A595857464544434241303F3E3D3C2B2A2928272;
defparam prom_inst_4.INIT_RAM_18 = 256'h6C5C4C3C2C1B0BFBEBDBCBBAAA9A8A7A6A594939291909F8E8D8C8B8A8978777;
defparam prom_inst_4.INIT_RAM_19 = 256'h7161514131201000F0E0D0C0AF9F8F7F6F5F4E3E2E1E0EFEEEDDCDBDAD9D8D7C;
defparam prom_inst_4.INIT_RAM_1A = 256'h7666564635251505F5E5D4C4B4A494847463534333231303F2E2D2C2B2A29281;
defparam prom_inst_4.INIT_RAM_1B = 256'h7A6A5A4A3A2A1A09F9E9D9C9B9A998887868584838271707F7E7D7C7B6A69686;
defparam prom_inst_4.INIT_RAM_1C = 256'h7E6E5E4E3E2E1E0EFDEDDDCDBDAD9D8D7C6C5C4C3C2C1C0BFBEBDBCBBBAB9B8A;
defparam prom_inst_4.INIT_RAM_1D = 256'h827262524232211101F1E1D1C1B1A190807060504030200FFFEFDFCFBFAF9F8F;
defparam prom_inst_4.INIT_RAM_1E = 256'h867565554535251505F5E5D4C4B4A494847464544333231303F3E3D3C3B2A292;
defparam prom_inst_4.INIT_RAM_1F = 256'h897968584838281808F8E8D8C8B7A797877767574737271606F6E6D6C6B6A696;
defparam prom_inst_4.INIT_RAM_20 = 256'h8B7B6B5B4B3B2B1B0BFBEBDACABAAA9A8A7A6A5A4A3A2A1909F9E9D9C9B9A999;
defparam prom_inst_4.INIT_RAM_21 = 256'h8E7E6E5E4D3D2D1D0DFDEDDDCDBDAD9D8D7D6C5C4C3C2C1C0CFCECDCCCBCAC9B;
defparam prom_inst_4.INIT_RAM_22 = 256'h90807060503F2F1F0FFFEFDFCFBFAF9F8F7F6F5F4F3F2E1E0EFEEEDECEBEAE9E;
defparam prom_inst_4.INIT_RAM_23 = 256'h91817161514131211101F1E1D1C1B1A191817160504030201000F0E0D0C0B0A0;
defparam prom_inst_4.INIT_RAM_24 = 256'h93837363534232221202F2E2D2C2B2A292827262524232221202F2E2D2C2B2A1;
defparam prom_inst_4.INIT_RAM_25 = 256'h94847363534333231303F3E3D3C3B3A393837363534333231303F3E3D3C3B3A3;
defparam prom_inst_4.INIT_RAM_26 = 256'h94847464544434241404F4E4D4C4B4A494847464544434241404F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_27 = 256'h94847464544434241404F4E4D4C4B4A494847464544434241404F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_28 = 256'h94847464544434241404F4E4D4C4B4A494847464544434241404F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_29 = 256'h93837363534333231303F3E3D3C3B3A393837363534333231304F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_2A = 256'h92827262524232221202F2E2D2C2B2A292827262524233231303F3E3D3C3B3A3;
defparam prom_inst_4.INIT_RAM_2B = 256'h90807060504030201000F0E1D1C1B1A191817161514131211101F1E1D1C1B2A2;
defparam prom_inst_4.INIT_RAM_2C = 256'h8E7E6E5E4E3E2E1E0EFEEEDFCFBFAF9F8F7F6F5F4F3F2F1F0FFFF0E0D0C0B0A0;
defparam prom_inst_4.INIT_RAM_2D = 256'h8B7B6B5B4C3C2C1C0CFCECDCCCBCAC9C8D7D6D5D4D3D2D1D0DFDEDDDCDBEAE9E;
defparam prom_inst_4.INIT_RAM_2E = 256'h887868584839291909F9E9D9C9B9A99A8A7A6A5A4A3A2A1A0AFBEBDBCBBBAB9B;
defparam prom_inst_4.INIT_RAM_2F = 256'h857565554535251505F6E6D6C6B6A696867667574737271707F7E7D8C8B8A898;
defparam prom_inst_4.INIT_RAM_30 = 256'h807161514131211102F2E2D2C2B2A292837363534333231304F4E4D4C4B4A494;
defparam prom_inst_4.INIT_RAM_31 = 256'h7C6C5C4C3C2D1D0DFDEDDDCEBEAE9E8E7E6E5F4F3F2F1F0FFFF0E0D0C0B0A090;
defparam prom_inst_4.INIT_RAM_32 = 256'h7767574737281808F8E8D8C9B9A99989796A5A4A3A2A1A0BFBEBDBCBBBAB9C8C;
defparam prom_inst_4.INIT_RAM_33 = 256'h7161524232221203F3E3D3C3B3A494847464544535251505F5E6D6C6B6A69687;
defparam prom_inst_4.INIT_RAM_34 = 256'h6B5B4C3C2C1C0CFDEDDDCDBDAD9E8E7E6E5E4F3F2F1F0F00F0E0D0C0B0A19181;
defparam prom_inst_4.INIT_RAM_35 = 256'h64554535251606F6E6D6C7B7A797877868584838291909F9EADACABAAA9B8B7B;
defparam prom_inst_4.INIT_RAM_36 = 256'h5D4E3E2E1E0EFFEFDFCFC0B0A090807161514132221202F2E3D3C3B3A4948474;
defparam prom_inst_4.INIT_RAM_37 = 256'h564636261707F7E7D8C8B8A898897969594A3A2A1A0BFBEBDBCCBCAC9C8D7D6D;
defparam prom_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000E3D3C4B4A495857565;
defparam prom_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[23:0],dout[47:40]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 8;
defparam prom_inst_5.RESET_MODE = "ASYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0C0C0C0C0C;
defparam prom_inst_5.INIT_RAM_01 = 256'h1010101010101010101010100F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0E0E0E0E;
defparam prom_inst_5.INIT_RAM_02 = 256'h1212121212121212121212121211111111111111111111111111111110101010;
defparam prom_inst_5.INIT_RAM_03 = 256'h1414141414141414141414141413131313131313131313131313131313121212;
defparam prom_inst_5.INIT_RAM_04 = 256'h1616161616161616161616161616151515151515151515151515151515151414;
defparam prom_inst_5.INIT_RAM_05 = 256'h1818181818181818181818181818171717171717171717171717171717171616;
defparam prom_inst_5.INIT_RAM_06 = 256'h1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1919191919191919191919191919191918;
defparam prom_inst_5.INIT_RAM_07 = 256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1A;
defparam prom_inst_5.INIT_RAM_08 = 256'h1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D;
defparam prom_inst_5.INIT_RAM_09 = 256'h21202020202020202020202020202020201F1F1F1F1F1F1F1F1F1F1F1F1F1F1F;
defparam prom_inst_5.INIT_RAM_0A = 256'h2322222222222222222222222222222222212121212121212121212121212121;
defparam prom_inst_5.INIT_RAM_0B = 256'h2525242424242424242424242424242424242323232323232323232323232323;
defparam prom_inst_5.INIT_RAM_0C = 256'h2727262626262626262626262626262626262525252525252525252525252525;
defparam prom_inst_5.INIT_RAM_0D = 256'h2929292828282828282828282828282828282827272727272727272727272727;
defparam prom_inst_5.INIT_RAM_0E = 256'h2B2B2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A29292929292929292929292929;
defparam prom_inst_5.INIT_RAM_0F = 256'h2D2D2D2D2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2B2B2B2B2B;
defparam prom_inst_5.INIT_RAM_10 = 256'h2F2F2F2F2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2D2D2D2D2D2D2D2D2D2D2D2D;
defparam prom_inst_5.INIT_RAM_11 = 256'h31313131313030303030303030303030303030302F2F2F2F2F2F2F2F2F2F2F2F;
defparam prom_inst_5.INIT_RAM_12 = 256'h3333333333323232323232323232323232323232323131313131313131313131;
defparam prom_inst_5.INIT_RAM_13 = 256'h3535353535343434343434343434343434343434343333333333333333333333;
defparam prom_inst_5.INIT_RAM_14 = 256'h3737373737373636363636363636363636363636363635353535353535353535;
defparam prom_inst_5.INIT_RAM_15 = 256'h3939393939393838383838383838383838383838383837373737373737373737;
defparam prom_inst_5.INIT_RAM_16 = 256'h3B3B3B3B3B3B3B3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A39393939393939393939;
defparam prom_inst_5.INIT_RAM_17 = 256'h3D3D3D3D3D3D3D3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3B3B3B3B3B3B3B3B3B;
defparam prom_inst_5.INIT_RAM_18 = 256'h3F3F3F3F3F3F3F3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3D3D3D3D3D3D3D3D3D;
defparam prom_inst_5.INIT_RAM_19 = 256'h41414141414141414040404040404040404040404040403F3F3F3F3F3F3F3F3F;
defparam prom_inst_5.INIT_RAM_1A = 256'h4343434343434343424242424242424242424242424242424141414141414141;
defparam prom_inst_5.INIT_RAM_1B = 256'h4545454545454545444444444444444444444444444444444343434343434343;
defparam prom_inst_5.INIT_RAM_1C = 256'h4747474747474747464646464646464646464646464646464545454545454545;
defparam prom_inst_5.INIT_RAM_1D = 256'h4949494949494949494848484848484848484848484848484747474747474747;
defparam prom_inst_5.INIT_RAM_1E = 256'h4B4B4B4B4B4B4B4B4B4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A49494949494949;
defparam prom_inst_5.INIT_RAM_1F = 256'h4D4D4D4D4D4D4D4D4D4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4B4B4B4B4B4B4B;
defparam prom_inst_5.INIT_RAM_20 = 256'h4F4F4F4F4F4F4F4F4F4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4D4D4D4D4D4D4D;
defparam prom_inst_5.INIT_RAM_21 = 256'h515151515151515151505050505050505050505050505050504F4F4F4F4F4F4F;
defparam prom_inst_5.INIT_RAM_22 = 256'h5353535353535353535252525252525252525252525252525251515151515151;
defparam prom_inst_5.INIT_RAM_23 = 256'h5555555555555555555554545454545454545454545454545454535353535353;
defparam prom_inst_5.INIT_RAM_24 = 256'h5757575757575757575756565656565656565656565656565656555555555555;
defparam prom_inst_5.INIT_RAM_25 = 256'h5959595959595959595958585858585858585858585858585858575757575757;
defparam prom_inst_5.INIT_RAM_26 = 256'h5B5B5B5B5B5B5B5B5B5B5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A595959595959;
defparam prom_inst_5.INIT_RAM_27 = 256'h5D5D5D5D5D5D5D5D5D5D5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5B5B5B5B5B5B;
defparam prom_inst_5.INIT_RAM_28 = 256'h5F5F5F5F5F5F5F5F5F5F5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5D5D5D5D5D5D;
defparam prom_inst_5.INIT_RAM_29 = 256'h61616161616161616161606060606060606060606060606060605F5F5F5F5F5F;
defparam prom_inst_5.INIT_RAM_2A = 256'h6363636363636363636362626262626262626262626262626262616161616161;
defparam prom_inst_5.INIT_RAM_2B = 256'h6565656565656565656564646464646464646464646464646464636363636363;
defparam prom_inst_5.INIT_RAM_2C = 256'h6767676767676767676666666666666666666666666666666665656565656565;
defparam prom_inst_5.INIT_RAM_2D = 256'h6969696969696969696868686868686868686868686868686867676767676767;
defparam prom_inst_5.INIT_RAM_2E = 256'h6B6B6B6B6B6B6B6B6B6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A69696969696969;
defparam prom_inst_5.INIT_RAM_2F = 256'h6D6D6D6D6D6D6D6D6D6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6B6B6B6B6B6B6B;
defparam prom_inst_5.INIT_RAM_30 = 256'h6F6F6F6F6F6F6F6F6F6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6D6D6D6D6D6D6D;
defparam prom_inst_5.INIT_RAM_31 = 256'h7171717171717171707070707070707070707070707070706F6F6F6F6F6F6F6F;
defparam prom_inst_5.INIT_RAM_32 = 256'h7373737373737373727272727272727272727272727272727171717171717171;
defparam prom_inst_5.INIT_RAM_33 = 256'h7575757575757575747474747474747474747474747474747373737373737373;
defparam prom_inst_5.INIT_RAM_34 = 256'h7777777777777776767676767676767676767676767676767575757575757575;
defparam prom_inst_5.INIT_RAM_35 = 256'h7979797979797978787878787878787878787878787878777777777777777777;
defparam prom_inst_5.INIT_RAM_36 = 256'h7B7B7B7B7B7B7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A797979797979797979;
defparam prom_inst_5.INIT_RAM_37 = 256'h7D7D7D7D7D7D7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7B7B7B7B7B7B7B7B7B7B;
defparam prom_inst_5.INIT_RAM_38 = 256'h00000000000000000000000000000000000000000000007D7D7D7D7D7D7D7D7D;
defparam prom_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //romcoef_module

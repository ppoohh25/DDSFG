//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10 (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Wed Jul 31 20:16:20 2024

module romcoef_module (dout, clk, oce, ce, reset, ad);

output [47:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire [23:0] prom_inst_2_dout_w;
wire [23:0] prom_inst_3_dout_w;
wire [23:0] prom_inst_4_dout_w;
wire [23:0] prom_inst_5_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hAACEEE091F303D464A49443A2B1800E4C39E734511DA9D5C16CC7D29D17513AD;
defparam prom_inst_0.INIT_RAM_01 = 256'hAE6517C56F13B34FE678068F14940F86F866CF3393EE4597E42D71B1EC225482;
defparam prom_inst_0.INIT_RAM_02 = 256'h4E98DE1F5B93C6F51F44658299ACBBC5CACBC7BEB1A0896E4F2B02D5A36D31F2;
defparam prom_inst_0.INIT_RAM_03 = 256'h8C694216E5B07638F5AE6211BC6204A139CD5CE66CEE6BE356C53096F753ABFF;
defparam prom_inst_0.INIT_RAM_04 = 256'h68D844AB0D6BC51A6AB5FC3F7CB6EA1A466D8FACC5DAEAF5FCFEFBF4E8D8C3AA;
defparam prom_inst_0.INIT_RAM_05 = 256'hE3E6E5DFD5C6B29A7D5C360BDCA87033F1AB6011BD6508A640D565F178FB79F3;
defparam prom_inst_0.INIT_RAM_06 = 256'hFF9527B43CC040BA31A20F78DB3B95EB3D8AD215558FC5F6234B6E8DA8BDCFDB;
defparam prom_inst_0.INIT_RAM_07 = 256'hBBE5092A455C6E7C858A8A857C6E5B442909E4BA8C5A23E7A76218CA7720C464;
defparam prom_inst_0.INIT_RAM_08 = 256'h1BD78E41F09A3FE07C13A634BE43C33FB729980166C62279CC1A63A8E8245B8E;
defparam prom_inst_0.INIT_RAM_09 = 256'h1E6DB7FD3E7BB3E715406687A3BBCFDDE8EDEEEBE3D6C4AF94755129FCCB955A;
defparam prom_inst_0.INIT_RAM_0A = 256'hC5A7855D3101CC925411CA7E2DD87E20BD55E97803890B880074E34EB41572CA;
defparam prom_inst_0.INIT_RAM_0B = 256'h1388F864CB2D8BE43888D41A5D9AD308386389ACC9E2F60611181A171004F4DF;
defparam prom_inst_0.INIT_RAM_0C = 256'h091113120B00F1DDC4A7855E3304D0975917D18636E2892BC962F787139A1C9A;
defparam prom_inst_0.INIT_RAM_0D = 256'hA843D869F57D007FF96EDF4BB31674CE2474C0084B89C3F829557DA0BED8EDFD;
defparam prom_inst_0.INIT_RAM_0E = 256'hF31F476B8AA4BACBD8E0E3E2DDD2C3B0987B5A340ADBA87033F2AC6112BF670A;
defparam prom_inst_0.INIT_RAM_0F = 256'hE9A86319CB7820C463FE9425B23BBE3EB82EA00C75D83792E83986CE12518BC1;
defparam prom_inst_0.INIT_RAM_10 = 256'h8EE02D76BAFA356B9DCAF21636516779868E92928D8374624A2E0DE8BE905D25;
defparam prom_inst_0.INIT_RAM_11 = 256'hE4C8A883592BF9C2864501B76916BF63039E34C654DC61E05BD243B1197DDD38;
defparam prom_inst_0.INIT_RAM_12 = 256'hEC62D442AB0F6FCA2173C0094E8DC9FF315F88ACCCE7FD0F1D262A2A251C0EFB;
defparam prom_inst_0.INIT_RAM_13 = 256'hA8B1B5B5B0A799876F54340FE6B8854E13D38E45F7A44DF2922DC356E36CF070;
defparam prom_inst_0.INIT_RAM_14 = 256'h1AB54CDE6CF579F974EB5DCB3498F853AAFC4A93D7175289BBE912365671889A;
defparam prom_inst_0.INIT_RAM_15 = 256'h45729BC0DFFB1123313A3E3E3930220FF8DDBC986E400ED79B5B16CD7F2DD67A;
defparam prom_inst_0.INIT_RAM_16 = 256'h2BEBA65C0EBB6408A843D96BF98206850177E956BF2483DE3587D41D62A1DC13;
defparam prom_inst_0.INIT_RAM_17 = 256'hCE206DB5F93974AADC0931557590A6B8C5CDD1D1CCC2B4A18A6E4E29FFD19E67;
defparam prom_inst_0.INIT_RAM_18 = 256'h3115F4CEA476420BCE8E48FEB05C05A848E2780A971FA3229D1385F25ABE1D78;
defparam prom_inst_0.INIT_RAM_19 = 256'h57CC3DA91174D32D83D42068ACEA255A8BB8E003223D526470787C7B756B5C49;
defparam prom_inst_0.INIT_RAM_1A = 256'h41484B4943382814FBDEBD966C3C08D093510BC0711DC56806A036C753DB5EDC;
defparam prom_inst_0.INIT_RAM_1B = 256'hF28B20B03BC244C23BB0208BF255B20C60B1FC4386C4FD32628EB5D8F60F2435;
defparam prom_inst_0.INIT_RAM_1C = 256'h6E99BFE1FE162A39444A4C4942362610F7D9B68F6333FEC48644FDB1610CB355;
defparam prom_inst_0.INIT_RAM_1D = 256'hB8742BDF8D37DD7E1AB245D45EE465E159CD3CA60C6DCA2275C40F5596D30B3F;
defparam prom_inst_0.INIT_RAM_1E = 256'hD11F68ACEC285F91BFE80D2D496073818A8F8F8B8375644D3213EFC6996832F7;
defparam prom_inst_0.INIT_RAM_1F = 256'hBE9D774D1EEBB47736F1A75906AE52F28D23B542CB4FCF4AC032A0096DCD287F;
defparam prom_inst_0.INIT_RAM_20 = 256'h80F15CC42684DE3383CF175A98D20738648CAFCDE7FD0E1A2225241E1405F2DA;
defparam prom_inst_0.INIT_RAM_21 = 256'h1D1E1B1307F6E1C7A9865F3302CD945613CC8030DB8224C25BF0800B9214920C;
defparam prom_inst_0.INIT_RAM_22 = 256'h9628B640C445C138AB1983E848A4FC4F9DE72D6EAAE215446E94B5D2EAFD0C17;
defparam prom_inst_0.INIT_RAM_23 = 256'hEF12314C61737F888B8B857B6D5A432706E1B8895720E4A45F16C8751FC363FF;
defparam prom_inst_0.INIT_RAM_24 = 256'h2CE0903BE18421BA4FDF6AF174F26BE051BC2487E53F94E43178BBFA346A9BC7;
defparam prom_inst_0.INIT_RAM_25 = 256'h4F94D511487BA9D3F819364D616F797F807D75695842280AE7BF93622DF4B573;
defparam prom_inst_0.INIT_RAM_26 = 256'h5D3304D1995C1BD68C3DEA9236D671079926AF33B32EA51785EE52B20E65B806;
defparam prom_inst_0.INIT_RAM_27 = 256'h5AC0227FD72B7BC60C4E8CC5F929547B9EBCD5EAFA060D100E08FDEEDAC2A583;
defparam prom_inst_0.INIT_RAM_28 = 256'h493F311E07ECCCA77E501EE8AC6D29E09341EB9031CD65F887119718940D80EF;
defparam prom_inst_0.INIT_RAM_29 = 256'h2DB436B42DA2127DE547A5FF54A5F1397CBAF42A5B88B0D3F20D2335424A4E4E;
defparam prom_inst_0.INIT_RAM_2A = 256'h0B2234424C50514D4437250FF4D5B2895D2BF6BC7D3AF2A65500A648E57E12A2;
defparam prom_inst_0.INIT_RAM_2B = 256'hE78E30CE68FD8D19A023A11B91026ED63998F3489AE72F73B2ED245583ACD0F0;
defparam prom_inst_0.INIT_RAM_2C = 256'hC5FC2E5C85AACAE6FD101E282D2E2B221605EFD5B6936B3F0ED9A0611FD88C3C;
defparam prom_inst_0.INIT_RAM_2D = 256'hA97032EFA85D0DB85F02A03ACF5FEB73F675EF65D642AB0E6DC81E70BD064A8A;
defparam prom_inst_0.INIT_RAM_2E = 256'h97ED3F8CD5195994CBFD2B547999B5CCDFEDF7FCFDF9F1E5D4BEA485623B0FDE;
defparam prom_inst_0.INIT_RAM_2F = 256'h947A5B3710E3B27D4305C27B2FDF8A31D4710BA030BC44C745BF34A5127ADE3D;
defparam prom_inst_0.INIT_RAM_30 = 256'hA41989F55DC01E78CE1F6CB4F73771A8D9072F54748FA6B8C6D0D5D5D1C8BCAA;
defparam prom_inst_0.INIT_RAM_31 = 256'hCBCFCFCAC1B3A18A6F4F2B03D5A46E33F4B1691DCC761CBE5BF48818A32AAD2B;
defparam prom_inst_0.INIT_RAM_32 = 256'h0FA230BB40C23FB72B9A056CCE2B84D92975BCFF3D77ACDD093155748EA4B6C3;
defparam prom_inst_0.INIT_RAM_33 = 256'h7395B2CBE0F0FC030605FEF4E5D1B99D7C572DFFCC955919D48B3EEC953ADB77;
defparam prom_inst_0.INIT_RAM_34 = 256'hFCAD5901A544DE7406931CA0209B1284F25CC1217DD52877C1074885BEF1214C;
defparam prom_inst_0.INIT_RAM_35 = 256'hB0EF2A6193C0E90E2E4A6274838D929490887C6B563C1EFCD5A979450CCF8D47;
defparam prom_inst_0.INIT_RAM_36 = 256'h92602AEFAF6B23D6852FD57613AC40D05BE164E15BD040AC1477D52F85D6236C;
defparam prom_inst_0.INIT_RAM_37 = 256'hA9055DB0FF4A90D10E477BABD6FD1F3D576C7D899094938D8374614A2E0EE9C0;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000A327A723990C7AE348;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "ASYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h2024282D3135393D4145494D5155595C6064686C7073777B7F82868A8D919598;
defparam prom_inst_1.INIT_RAM_01 = 256'h92979CA0A5AAAEB3B7BCC1C5CACED3D7DBE0E4E9EDF1F6FAFE03070B0F14181C;
defparam prom_inst_1.INIT_RAM_02 = 256'hF2F7FC02070C11161C21262B30353A3F44494E53585D62676C71767A7F84898D;
defparam prom_inst_1.INIT_RAM_03 = 256'h3F454B51565C62686D73797F848A90959BA0A6ABB1B6BCC1C7CCD2D7DCE2E7EC;
defparam prom_inst_1.INIT_RAM_04 = 256'h7A80878D949AA0A7ADB3B9C0C6CCD2D9DFE5EBF1F7FD03090F151B21272D3339;
defparam prom_inst_1.INIT_RAM_05 = 256'hA2A9B0B7BEC5CCD3DAE1E8EFF5FC030A10171E252B32393F464C535960666D73;
defparam prom_inst_1.INIT_RAM_06 = 256'hB8C0C8CFD7DEE6EDF5FC040B121A212830373E464D545B626A71787F868D949B;
defparam prom_inst_1.INIT_RAM_07 = 256'hBCC4CDD5DDE5EDF5FD050D151D252D353D454C545C646C737B838B929AA2A9B1;
defparam prom_inst_1.INIT_RAM_08 = 256'hAEB6BFC8D0D9E2EAF3FC040D151E262F3740485159616A727A838B939BA4ACB4;
defparam prom_inst_1.INIT_RAM_09 = 256'h8D969FA8B2BBC4CDD7E0E9F2FB040D161F28313A434C555E677079828A939CA5;
defparam prom_inst_1.INIT_RAM_0A = 256'h59636D77818B949EA8B2BBC5CFD8E2ECF5FF08121C252F38424B545E67717A83;
defparam prom_inst_1.INIT_RAM_0B = 256'h141E28333D48525C67717B86909AA4AFB9C3CDD7E1EBF5000A141E28323C454F;
defparam prom_inst_1.INIT_RAM_0C = 256'hBCC7D2DDE8F3FD08131E29343F4A545F6A757F8A959FAAB5BFCAD4DFEAF4FF09;
defparam prom_inst_1.INIT_RAM_0D = 256'h515D68747F8B97A2ADB9C4D0DBE7F2FD09141F2B36414C57636E79848F9AA5B0;
defparam prom_inst_1.INIT_RAM_0E = 256'hD4E1EDF905111D2935414D5965717D8995A1ADB9C5D0DCE8F4FF0B17232E3A46;
defparam prom_inst_1.INIT_RAM_0F = 256'h45525F6C7885929EABB7C4D1DDEAF6030F1C2835414D5A66727F8B97A4B0BCC8;
defparam prom_inst_1.INIT_RAM_10 = 256'hA4B1BFCCD9E6F4010E1B283643505D6A7784919EABB8C5D2DFECF905121F2C39;
defparam prom_inst_1.INIT_RAM_11 = 256'hF0FE0C1A283643515F6D7B8896A4B1BFCDDAE8F503101E2B394654616F7C8997;
defparam prom_inst_1.INIT_RAM_12 = 256'h2A3947566473818F9EACBAC9D7E5F301101E2C3A48566473818F9DABB9C7D5E2;
defparam prom_inst_1.INIT_RAM_13 = 256'h5261707F8E9DACBBCAD9E8F705142332414F5E6D7B8A99A7B6C5D3E2F0FF0D1C;
defparam prom_inst_1.INIT_RAM_14 = 256'h68778796A6B5C5D4E4F30312223140505F6E7E8D9CACBBCAD9E8F80716253443;
defparam prom_inst_1.INIT_RAM_15 = 256'h6B7B8B9BABBBCCDCECFC0C1C2C3C4C5C6B7B8B9BABBBCBDAEAFA0A1929394858;
defparam prom_inst_1.INIT_RAM_16 = 256'h5C6C7D8E9FAFC0D1E1F202132334455566768697A7B8C8D8E9F9091A2A3A4A5B;
defparam prom_inst_1.INIT_RAM_17 = 256'h3A4C5D6E7F91A2B3C4D6E7F8091A2B3C4D5E6F8091A2B3C4D5E6F70818293A4B;
defparam prom_inst_1.INIT_RAM_18 = 256'h07192A3C4E60728495A7B9CADCEE001123344658697B8C9EAFC1D2E3F5061829;
defparam prom_inst_1.INIT_RAM_19 = 256'hC1D3E6F80B1D2F425466798B9DAFC2D4E6F80A1D2F41536577899BADBFD1E3F5;
defparam prom_inst_1.INIT_RAM_1A = 256'h697C8FA2B5C8DBEE001326394C5F728497AABDCFE2F5071A2D3F526477899CAE;
defparam prom_inst_1.INIT_RAM_1B = 256'hFE1226394D6074879BAEC2D5E8FC0F2336495C708396A9BDD0E3F6091C304356;
defparam prom_inst_1.INIT_RAM_1C = 256'h8296AABED2E7FB0F23374B5F73879BAFC2D6EAFE1226394D6175889CB0C4D7EB;
defparam prom_inst_1.INIT_RAM_1D = 256'hF3081D31465B6F8499ADC2D6EBFF14283D51667A8FA3B7CCE0F4091D31455A6E;
defparam prom_inst_1.INIT_RAM_1E = 256'h52687D92A7BDD2E7FC11273C51667B90A5BACFE4F90E23384D62768BA0B5CADE;
defparam prom_inst_1.INIT_RAM_1F = 256'h9FB5CBE1F70C22384E63798FA5BAD0E5FB11263C51677C92A7BDD2E8FD12283D;
defparam prom_inst_1.INIT_RAM_20 = 256'hDAF0071D344A60778DA3BAD0E6FC13293F556B8197ADC4DAF0061C32485E7389;
defparam prom_inst_1.INIT_RAM_21 = 256'h031A31485F758CA3BAD1E8FF162C435A71879EB5CBE2F90F263C536A8097ADC4;
defparam prom_inst_1.INIT_RAM_22 = 256'h19314860778FA6BED5ED041B334A617990A7BFD6ED041C334A61788FA6BDD5EC;
defparam prom_inst_1.INIT_RAM_23 = 256'h1D364E667E96AEC6DEF60E263E566E869EB5CDE5FD152C445C748BA3BBD2EA01;
defparam prom_inst_1.INIT_RAM_24 = 256'h1028415A728BA4BCD5ED061E374F688099B1CAE2FA132B435C748CA4BDD5ED05;
defparam prom_inst_1.INIT_RAM_25 = 256'hF009223C556E87A0B9D3EC051E375069829BB4CDE6FF183149627B94ADC5DEF7;
defparam prom_inst_1.INIT_RAM_26 = 256'hBED8F20B253F59728CA6BFD9F30C264059738CA6BFD9F20C253E58718BA4BDD7;
defparam prom_inst_1.INIT_RAM_27 = 256'h7A94AFC9E3FE18324D67819BB5D0EA041E38526C86A1BBD5EF09223C56708AA4;
defparam prom_inst_1.INIT_RAM_28 = 256'h243F5A7590AAC5E0FB16314B66819CB6D1EC06213C56718BA6C1DBF6102B455F;
defparam prom_inst_1.INIT_RAM_29 = 256'hBCD7F30E2A45617C97B3CEE905203B57728DA8C4DFFA15304B67829DB8D3EE09;
defparam prom_inst_1.INIT_RAM_2A = 256'h425E7A96B2CEEA06223E5A7691ADC9E5011D3854708CA7C3DFFB16324D6985A0;
defparam prom_inst_1.INIT_RAM_2B = 256'hB5D2EF0B2844617E9AB7D3F00C2945617E9AB6D3EF0B2844607C99B5D1ED0925;
defparam prom_inst_1.INIT_RAM_2C = 256'h1734526F8CA9C6E3001E3B587592AFCCE906223F5C7996B3D0EC0926435F7C99;
defparam prom_inst_1.INIT_RAM_2D = 256'h6785A3C0DEFC1A37557390AECBE90624415F7C9AB7D5F2102D4A6885A2C0DDFA;
defparam prom_inst_1.INIT_RAM_2E = 256'hA5C3E2001E3D5B7997B5D4F2102E4C6A88A6C4E2001E3C5A7896B4D2F00E2C49;
defparam prom_inst_1.INIT_RAM_2F = 256'hD1F00F2E4D6B8AA9C8E705244361809FBDDCFB1938567593B2D0EF0D2C4A6887;
defparam prom_inst_1.INIT_RAM_30 = 256'hEB0B2A496988A8C7E60625446383A2C1E0001F3E5D7C9BBAD9F81736557493B2;
defparam prom_inst_1.INIT_RAM_31 = 256'hF31333537393B3D3F31333537292B2D2F11131517090B0CFEF0E2E4E6D8DACCC;
defparam prom_inst_1.INIT_RAM_32 = 256'hEA0A2B4B6C8CADCDEE0E2F4F6F90B0D0F11131517292B2D2F31333537393B3D3;
defparam prom_inst_1.INIT_RAM_33 = 256'hCEEF1031527394B6D7F818395A7B9CBDDEFF20406182A3C4E40526466788A8C9;
defparam prom_inst_1.INIT_RAM_34 = 256'hA0C2E40627496A8CAECFF11234557798B9DBFC1E3F6082A3C4E60728496A8CAD;
defparam prom_inst_1.INIT_RAM_35 = 256'h6183A6C8EA0C2E517395B7D9FB1D3F6183A5C7E90B2D4F7092B4D6F81A3B5D7F;
defparam prom_inst_1.INIT_RAM_36 = 256'h103356789BBEE10326496B8EB1D3F6183B5D80A2C5E70A2C4F7193B6D8FA1D3F;
defparam prom_inst_1.INIT_RAM_37 = 256'hADD1F4173A5E81A4C8EB0E3154779BBEE104274A6D90B3D6F91C3F6285A8CAED;
defparam prom_inst_1.INIT_RAM_38 = 256'h00000000000000000000000000000000000000000000006E92B5D9FC2043668A;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[23:0],dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 8;
defparam prom_inst_2.RESET_MODE = "ASYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE;
defparam prom_inst_2.INIT_RAM_01 = 256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFEFEFEFEFEFEFE;
defparam prom_inst_2.INIT_RAM_02 = 256'hFCFCFCFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD;
defparam prom_inst_2.INIT_RAM_03 = 256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC;
defparam prom_inst_2.INIT_RAM_04 = 256'hFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFCFCFCFCFCFCFCFCFCFC;
defparam prom_inst_2.INIT_RAM_05 = 256'hFAFAFAFAFAFAFAFAFAFAFAFAFAFAFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB;
defparam prom_inst_2.INIT_RAM_06 = 256'hF9F9F9F9F9F9F9F9F9F9FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA;
defparam prom_inst_2.INIT_RAM_07 = 256'hF8F8F8F8F8F8F8F8F8F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9;
defparam prom_inst_2.INIT_RAM_08 = 256'hF7F7F7F7F7F7F7F7F7F7F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8;
defparam prom_inst_2.INIT_RAM_09 = 256'hF6F6F6F6F6F6F6F6F6F6F6F6F6F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7;
defparam prom_inst_2.INIT_RAM_0A = 256'hF5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F6F6F6F6F6F6F6F6F6F6F6F6F6F6;
defparam prom_inst_2.INIT_RAM_0B = 256'hF4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F5F5F5F5F5F5F5F5F5;
defparam prom_inst_2.INIT_RAM_0C = 256'hF2F2F2F2F2F2F2F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F4;
defparam prom_inst_2.INIT_RAM_0D = 256'hF1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2;
defparam prom_inst_2.INIT_RAM_0E = 256'hEFEFEFEFF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F1F1F1F1F1F1;
defparam prom_inst_2.INIT_RAM_0F = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF;
defparam prom_inst_2.INIT_RAM_10 = 256'hECECECECECECECEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_11 = 256'hEAEAEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBECECECECECECECECECECECEC;
defparam prom_inst_2.INIT_RAM_12 = 256'hE9E9E9E9E9E9E9E9E9E9E9E9E9E9E9EAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEA;
defparam prom_inst_2.INIT_RAM_13 = 256'hE7E7E7E7E7E7E7E7E7E7E7E7E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E9E9;
defparam prom_inst_2.INIT_RAM_14 = 256'hE5E5E5E5E5E5E5E5E5E5E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E7E7E7E7E7;
defparam prom_inst_2.INIT_RAM_15 = 256'hE3E3E3E3E3E3E3E3E3E3E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E5E5E5E5E5E5;
defparam prom_inst_2.INIT_RAM_16 = 256'hE1E1E1E1E1E1E1E1E1E1E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E3E3E3E3E3E3;
defparam prom_inst_2.INIT_RAM_17 = 256'hDFDFDFDFDFDFDFDFDFDFDFDFE0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E1E1E1E1E1;
defparam prom_inst_2.INIT_RAM_18 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDFDFDF;
defparam prom_inst_2.INIT_RAM_19 = 256'hDADADADADBDBDBDBDBDBDBDBDBDBDBDBDBDBDCDCDCDCDCDCDCDCDCDCDCDCDCDC;
defparam prom_inst_2.INIT_RAM_1A = 256'hD8D8D8D8D8D8D8D8D9D9D9D9D9D9D9D9D9D9D9D9D9D9DADADADADADADADADADA;
defparam prom_inst_2.INIT_RAM_1B = 256'hD5D6D6D6D6D6D6D6D6D6D6D6D6D6D7D7D7D7D7D7D7D7D7D7D7D7D7D8D8D8D8D8;
defparam prom_inst_2.INIT_RAM_1C = 256'hD3D3D3D3D3D3D3D4D4D4D4D4D4D4D4D4D4D4D4D4D5D5D5D5D5D5D5D5D5D5D5D5;
defparam prom_inst_2.INIT_RAM_1D = 256'hD0D1D1D1D1D1D1D1D1D1D1D1D1D1D2D2D2D2D2D2D2D2D2D2D2D2D3D3D3D3D3D3;
defparam prom_inst_2.INIT_RAM_1E = 256'hCECECECECECECECECECFCFCFCFCFCFCFCFCFCFCFCFD0D0D0D0D0D0D0D0D0D0D0;
defparam prom_inst_2.INIT_RAM_1F = 256'hCBCBCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCDCDCDCDCDCDCDCDCDCDCDCDCECECE;
defparam prom_inst_2.INIT_RAM_20 = 256'hC8C8C9C9C9C9C9C9C9C9C9C9C9C9CACACACACACACACACACACACBCBCBCBCBCBCB;
defparam prom_inst_2.INIT_RAM_21 = 256'hC6C6C6C6C6C6C6C6C6C6C6C6C7C7C7C7C7C7C7C7C7C7C7C8C8C8C8C8C8C8C8C8;
defparam prom_inst_2.INIT_RAM_22 = 256'hC3C3C3C3C3C3C3C3C3C3C4C4C4C4C4C4C4C4C4C4C4C5C5C5C5C5C5C5C5C5C5C5;
defparam prom_inst_2.INIT_RAM_23 = 256'hC0C0C0C0C0C0C0C0C0C0C1C1C1C1C1C1C1C1C1C1C1C2C2C2C2C2C2C2C2C2C2C3;
defparam prom_inst_2.INIT_RAM_24 = 256'hBDBDBDBDBDBDBDBDBDBDBEBEBEBEBEBEBEBEBEBEBEBFBFBFBFBFBFBFBFBFBFC0;
defparam prom_inst_2.INIT_RAM_25 = 256'hB9BABABABABABABABABABABBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBCBCBCBCBCBC;
defparam prom_inst_2.INIT_RAM_26 = 256'hB6B6B6B7B7B7B7B7B7B7B7B7B7B8B8B8B8B8B8B8B8B8B8B9B9B9B9B9B9B9B9B9;
defparam prom_inst_2.INIT_RAM_27 = 256'hB3B3B3B3B3B3B4B4B4B4B4B4B4B4B4B5B5B5B5B5B5B5B5B5B5B6B6B6B6B6B6B6;
defparam prom_inst_2.INIT_RAM_28 = 256'hB0B0B0B0B0B0B0B0B0B1B1B1B1B1B1B1B1B1B2B2B2B2B2B2B2B2B2B2B3B3B3B3;
defparam prom_inst_2.INIT_RAM_29 = 256'hACACACADADADADADADADADADAEAEAEAEAEAEAEAEAEAEAFAFAFAFAFAFAFAFAFB0;
defparam prom_inst_2.INIT_RAM_2A = 256'hA9A9A9A9A9A9A9AAAAAAAAAAAAAAAAAAABABABABABABABABABABACACACACACAC;
defparam prom_inst_2.INIT_RAM_2B = 256'hA5A5A5A6A6A6A6A6A6A6A6A6A7A7A7A7A7A7A7A7A7A8A8A8A8A8A8A8A8A8A9A9;
defparam prom_inst_2.INIT_RAM_2C = 256'hA2A2A2A2A2A2A2A2A3A3A3A3A3A3A3A3A3A4A4A4A4A4A4A4A4A4A5A5A5A5A5A5;
defparam prom_inst_2.INIT_RAM_2D = 256'h9E9E9E9E9E9E9F9F9F9F9F9F9F9FA0A0A0A0A0A0A0A0A0A1A1A1A1A1A1A1A1A1;
defparam prom_inst_2.INIT_RAM_2E = 256'h9A9A9A9B9B9B9B9B9B9B9B9B9C9C9C9C9C9C9C9C9D9D9D9D9D9D9D9D9D9E9E9E;
defparam prom_inst_2.INIT_RAM_2F = 256'h9696979797979797979798989898989898989899999999999999999A9A9A9A9A;
defparam prom_inst_2.INIT_RAM_30 = 256'h9293939393939393939494949494949494959595959595959595969696969696;
defparam prom_inst_2.INIT_RAM_31 = 256'h8E8F8F8F8F8F8F8F8F9090909090909090919191919191919192929292929292;
defparam prom_inst_2.INIT_RAM_32 = 256'h8A8B8B8B8B8B8B8B8B8C8C8C8C8C8C8C8C8D8D8D8D8D8D8D8D8E8E8E8E8E8E8E;
defparam prom_inst_2.INIT_RAM_33 = 256'h868687878787878787878888888888888888898989898989898A8A8A8A8A8A8A;
defparam prom_inst_2.INIT_RAM_34 = 256'h8282828383838383838383848484848484848485858585858585868686868686;
defparam prom_inst_2.INIT_RAM_35 = 256'h7E7E7E7E7E7F7F7F7F7F7F7F7F80808080808080818181818181818182828282;
defparam prom_inst_2.INIT_RAM_36 = 256'h7A7A7A7A7A7A7A7B7B7B7B7B7B7B7B7C7C7C7C7C7C7C7D7D7D7D7D7D7D7D7E7E;
defparam prom_inst_2.INIT_RAM_37 = 256'h7575757676767676767677777777777777787878787878787879797979797979;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000747474747475757575;
defparam prom_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[23:0],dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 8;
defparam prom_inst_3.RESET_MODE = "ASYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h974C02B76C21D68C41F6AB6015CA7F34E99E5308BD7227DC9146FAAF6419CE83;
defparam prom_inst_3.INIT_RAM_01 = 256'hE69C5208BD7329DE944AFFB56B20D68B41F6AC6117CC8237EDA2570DC2772DE2;
defparam prom_inst_3.INIT_RAM_02 = 256'h22D88F45FCB2681FD58B41F8AE641AD0873DF3A95F15CB8137EDA3590FC57A30;
defparam prom_inst_3.INIT_RAM_03 = 256'h48FFB66D24DC934A01B86F25DC934A01B86F25DC934A00B76E24DB9148FEB56B;
defparam prom_inst_3.INIT_RAM_04 = 256'h560EC67E36EEA55D15CD843CF4AB631BD28A41F9B0681FD78E45FDB46B22DA91;
defparam prom_inst_3.INIT_RAM_05 = 256'h4A03BC742DE69E5710C88139F2AA631BD48C44FDB56D25DE964E06BE762EE69E;
defparam prom_inst_3.INIT_RAM_06 = 256'h21DB954F08C27B35EEA8611BD48E4700B9732CE59E5711CA833CF5AE6720D891;
defparam prom_inst_3.INIT_RAM_07 = 256'hDA944F0AC47F3AF4AF6924DE98530DC7823CF6B06A24DE98520CC6803AF4AE68;
defparam prom_inst_3.INIT_RAM_08 = 256'h712DE8A4601CD7934E0AC5813CF8B36E2AE5A05B16D28D4803BE7934EFA9641F;
defparam prom_inst_3.INIT_RAM_09 = 256'hE4A15E1BD895510ECB884401BD7A36F3AF6C28E4A05D19D5914D09C5813DF9B5;
defparam prom_inst_3.INIT_RAM_0A = 256'h32F0AE6C2AE8A66422E09E5C19D7955210CD8B4806C3813EFBB97633F0AD6A27;
defparam prom_inst_3.INIT_RAM_0B = 256'h5716D6955514D3925111D08F4E0DCC8B4908C7864403C2803FFDBC7A39F7B573;
defparam prom_inst_3.INIT_RAM_0C = 256'h5112D3945415D6965717D8985919D9995A1ADA9A5A1ADA9A5A19D9995918D897;
defparam prom_inst_3.INIT_RAM_0D = 256'h1FE1A36628EAAC6E30F2B47537F9BB7C3EFFC1824405C788490ACB8D4E0FD090;
defparam prom_inst_3.INIT_RAM_0E = 256'hBD814508CC905317DA9E6124E7AB6E31F4B77A3D00C386480BCE905315D89A5D;
defparam prom_inst_3.INIT_RAM_0F = 256'h2AEFB47A3F04C98E5318DDA2672CF0B57A3E03C78C5015D99D6125E9AD7135F9;
defparam prom_inst_3.INIT_RAM_10 = 256'h6229F0B77E450CD2996026EDB37A4006CD93591FE5AB7137FDC3884E14D99F64;
defparam prom_inst_3.INIT_RAM_11 = 256'h652DF6BF875018E1A9723A02CA925A22EAB27A420AD1996128F0B77E460DD49B;
defparam prom_inst_3.INIT_RAM_12 = 256'h2EF9C38E5823EDB7814B15DFA9733D07D19A642DF7C08A531CE6AF78410AD39C;
defparam prom_inst_3.INIT_RAM_13 = 256'hBD895622EEBB87531FEBB7834E1AE6B27D4914DFAB76410CD8A36E3803CE9964;
defparam prom_inst_3.INIT_RAM_14 = 256'h0EDDAB794816E4B2804E1CE9B7855220EDBB885523F0BD8A5724F1BE8A5724F0;
defparam prom_inst_3.INIT_RAM_15 = 256'h20F0C191613202D2A2724111E1B180501FEFBE8D5D2CFBCA99683705D4A37140;
defparam prom_inst_3.INIT_RAM_16 = 256'hF0C295673A0CDEB0825426F8CA9B6D3F10E2B3855627F8C99A6B3C0DDEAE7F50;
defparam prom_inst_3.INIT_RAM_17 = 256'h7B5025F9CEA2764B1FF3C79B6F4317EBBE9265390CE0B386592CFFD2A5784B1D;
defparam prom_inst_3.INIT_RAM_18 = 256'hC0976E451CF2C99F764C22F9CFA57B5127FDD2A87E5329FED3A87E5328FDD2A7;
defparam prom_inst_3.INIT_RAM_19 = 256'hBC956F4821FAD3AB845D350EE6BF976F471FF8CFA77F572F06DEB58C643B12E9;
defparam prom_inst_3.INIT_RAM_1A = 256'h6D482400DBB6926D4823FED9B48E69441EF8D3AD87613C16EFC9A37D563009E3;
defparam prom_inst_3.INIT_RAM_1B = 256'hD0AE8C6A482603E1BF9C79573411EECBA885623F1BF8D4B18D694521FED9B591;
defparam prom_inst_3.INIT_RAM_1C = 256'hE3C4A48565462606E6C6A68665452504E4C3A28261401FFEDCBB9A78573514F2;
defparam prom_inst_3.INIT_RAM_1D = 256'hA4876B4E3114F6D9BC9E816346280AECCEB09274553718FADBBD9E7F60412202;
defparam prom_inst_3.INIT_RAM_1E = 256'h11F7DCC2A88D73583E2308EDD2B79C81654A2E13F7DBBFA3876B4F3316FADDC1;
defparam prom_inst_3.INIT_RAM_1F = 256'h260FF8E0C8B199816951392109F0D8BFA78E755C432A11F8DEC5AB92785E452B;
defparam prom_inst_3.INIT_RAM_20 = 256'hE3CEBAA5907B66513C2712FCE7D1BBA6907A644E38210BF4DEC7B19A836C553E;
defparam prom_inst_3.INIT_RAM_21 = 256'h4432210FFDEBD9C7B4A2907D6A5845321F0CF9E5D2BFAB9784705C4834200CF7;
defparam prom_inst_3.INIT_RAM_22 = 256'h47382A1B0CFDEEDFCFC0B0A191817161514131211000EFDECEBDAC9B89786755;
defparam prom_inst_3.INIT_RAM_23 = 256'hEADFD3C7BBAFA3978B7E7265584C3F3225180AFDF0E2D5C7B9AB9D8F81736456;
defparam prom_inst_3.INIT_RAM_24 = 256'h2B231A1108FFF6EDE4DBD1C8BEB5ABA1978D83796E64594F44392E23180D01F6;
defparam prom_inst_3.INIT_RAM_25 = 256'h0702FCF7F1EBE6E0DAD3CDC7C0BAB3ADA69F989189827B736C645C544C443C33;
defparam prom_inst_3.INIT_RAM_26 = 256'h7C7A787673716E6B696663605C5956524F4B47433F3B37322E2A25201B16110C;
defparam prom_inst_3.INIT_RAM_27 = 256'h88898A8B8C8D8E8E8F8F9090909090908F8F8E8E8D8C8B8A898886858382807E;
defparam prom_inst_3.INIT_RAM_28 = 256'h282D31363A3E42464A4E5255595C5F6266686B6E717376787A7C7E8082838587;
defparam prom_inst_3.INIT_RAM_29 = 256'h5A626A727A828991989FA6ADB4BBC2C9CFD5DCE2E8EEF4F9FF040A0F14191E23;
defparam prom_inst_3.INIT_RAM_2A = 256'h1C28333F4A55616C76818C96A1ABB5BFC9D3DDE7F0FA030C151E273039414A52;
defparam prom_inst_3.INIT_RAM_2B = 256'h6C7B8A99A8B7C6D4E3F1FF0E1C29374552606D7B8895A2AEBBC8D4E0EDF90510;
defparam prom_inst_3.INIT_RAM_2C = 256'h47596C7F92A4B7C9DBEDFF112234455768798A9BACBCCDDDEEFE0E1E2E3D4D5C;
defparam prom_inst_3.INIT_RAM_2D = 256'hAAC1D8EE041B31475D72889EB3C8DDF2071C31465A6E8397ABBFD2E6FA0D2033;
defparam prom_inst_3.INIT_RAM_2E = 256'h95AFC9E4FE18324C657F98B2CBE4FD162F47607890A9C1D8F0081F374E657C93;
defparam prom_inst_3.INIT_RAM_2F = 256'h0322405E7C9AB8D6F3112E4B6885A2BFDBF814304D6984A0BCD7F30E29445F7A;
defparam prom_inst_3.INIT_RAM_30 = 256'hF416395B7D9FC0E20425466789A9CAEB0B2C4C6C8CACCCEC0B2B4A6988A7C6E5;
defparam prom_inst_3.INIT_RAM_31 = 256'h648BB1D7FD23496F94BADF04294E7398BCE105294D7195B9DC002346698CAFD1;
defparam prom_inst_3.INIT_RAM_32 = 256'h527DA7D2FC26507AA3CDF61F49729AC3EC143D658DB5DD052C547BA2C9F0173E;
defparam prom_inst_3.INIT_RAM_33 = 256'hBCEA194776A4D2002E5C89B7E4113E6B98C4F11D4A76A2CDF925507CA7D2FD28;
defparam prom_inst_3.INIT_RAM_34 = 256'h9ED10436699BCE00326496C7F92A5C8DBEEF1F5080B1E1114171A0D0FF2F5E8D;
defparam prom_inst_3.INIT_RAM_35 = 256'hF72E659CD30A4177ADE41A5086BBF1265C91C6FB2F6498CD0135699DD004376B;
defparam prom_inst_3.INIT_RAM_36 = 256'hC4003B77B2ED28639ED8134D87C1FB356FA8E21B548DC6FF3770A8E0185088BF;
defparam prom_inst_3.INIT_RAM_37 = 256'h034484C3034382C201407FBEFC3B79B7F53371AFEC2A67A4E11E5B97D4104C88;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000BBFD3E7FC0014283C3;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[23:0],dout[39:32]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 8;
defparam prom_inst_4.RESET_MODE = "ASYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hB4A494837363524232211101F1E0D0C0AF9F8F7F6E5E4E3D2D1D0CFCECDCCBBB;
defparam prom_inst_4.INIT_RAM_01 = 256'hBDAD9D8D7C6C5C4B3B2B1A0AFAEAD9C9B9A898887867574736261606F5E5D5C4;
defparam prom_inst_4.INIT_RAM_02 = 256'hC7B6A696857565554434241303F3E3D2C2B2A19181716050402F1F0FFFEEDECE;
defparam prom_inst_4.INIT_RAM_03 = 256'hD0BFAF9F8F7E6E5E4E3D2D1D0CFCECDCCBBBAB9A8A7A6A594939281808F7E7D7;
defparam prom_inst_4.INIT_RAM_04 = 256'hD9C9B8A898877767574636261505F5E5D4C4B4A393837362524231211101F0E0;
defparam prom_inst_4.INIT_RAM_05 = 256'hE2D2C1B1A1908070604F3F2F1E0EFEEEDDCDBDAC9C8C7C6B5B4B3B2A1A0AF9E9;
defparam prom_inst_4.INIT_RAM_06 = 256'hEBDACABAAA99897968584838271707F7E6D6C6B5A595857464544333231302F2;
defparam prom_inst_4.INIT_RAM_07 = 256'hF3E3D3C3B2A2928171615140302010FFEFDFCEBEAE9E8D7D6D5D4C3C2C1B0BFB;
defparam prom_inst_4.INIT_RAM_08 = 256'hFCECDBCBBBAB9A8A7A6A594939281808F8E7D7C7B7A696867665554534241404;
defparam prom_inst_4.INIT_RAM_09 = 256'h04F4E4D4C3B3A393827262524131211000F0E0CFBFAF9F8E7E6E5E4D3D2D1C0C;
defparam prom_inst_4.INIT_RAM_0A = 256'h0DFCECDCCCBBAB9B8B7A6A5A4A39291909F8E8D8C8B7A7978676665645352515;
defparam prom_inst_4.INIT_RAM_0B = 256'h1505F4E4D4C4B3A393837262524231211101F0E0D0C0AF9F8F7E6E5E4E3D2D1D;
defparam prom_inst_4.INIT_RAM_0C = 256'h1D0DFCECDCCCBBAB9B8B7A6A5A4A39291909F8E8D8C8B7A79787766656463525;
defparam prom_inst_4.INIT_RAM_0D = 256'h251404F4E4D3C3B3A392827262514131211000F0E0D0BFAF9F8F7E6E5E4E3D2D;
defparam prom_inst_4.INIT_RAM_0E = 256'h2C1C0CFCEBDBCBBBAA9A8A7A69594939281808F8E8D7C7B7A796867666554535;
defparam prom_inst_4.INIT_RAM_0F = 256'h34231303F3E3D2C2B2A2918171615040302010FFEFDFCFBEAE9E8E7D6D5D4D3C;
defparam prom_inst_4.INIT_RAM_10 = 256'h3B2B1A0AFAEADAC9B9A999887868584837271707F6E6D6C6B5A5958575645444;
defparam prom_inst_4.INIT_RAM_11 = 256'h4232211101F1E1D0C0B0A0907F6F5F4F3E2E1E0EFEEDDDCDBDAC9C8C7C6C5B4B;
defparam prom_inst_4.INIT_RAM_12 = 256'h4938281808F8E7D7C7B7A796867666564535251504F4E4D4C4B3A39383736252;
defparam prom_inst_4.INIT_RAM_13 = 256'h4F3F2F1F0EFEEEDECEBDAD9D8D7D6C5C4C3C2C1B0BFBEBDBCABAAA9A8A796959;
defparam prom_inst_4.INIT_RAM_14 = 256'h564535251505F4E4D4C4B4A393837363524232221201F1E1D1C1B0A09080705F;
defparam prom_inst_4.INIT_RAM_15 = 256'h5C4B3B2B1B0BFBEADACABAAA99897969594838281808F7E7D7C7B7A796867666;
defparam prom_inst_4.INIT_RAM_16 = 256'h61514131211100F0E0D0C0AF9F8F7F6F5F4E3E2E1E0EFDEDDDCDBDAD9C8C7C6C;
defparam prom_inst_4.INIT_RAM_17 = 256'h67574736261606F6E6D5C5B5A595857464544434241303F3E3D3C2B2A2928272;
defparam prom_inst_4.INIT_RAM_18 = 256'h6C5C4C3C2C1B0BFBEBDBCBBAAA9A8A7A6A594939291909F8E8D8C8B8A8978777;
defparam prom_inst_4.INIT_RAM_19 = 256'h7161514131201000F0E0D0C0AF9F8F7F6F5F4E3E2E1E0EFEEEDDCDBDAD9D8D7C;
defparam prom_inst_4.INIT_RAM_1A = 256'h7666564635251505F5E5D4C4B4A494847463534333231303F2E2D2C2B2A29281;
defparam prom_inst_4.INIT_RAM_1B = 256'h7A6A5A4A3A2A1A09F9E9D9C9B9A998887868584838271707F7E7D7C7B6A69686;
defparam prom_inst_4.INIT_RAM_1C = 256'h7E6E5E4E3E2E1E0EFDEDDDCDBDAD9D8D7C6C5C4C3C2C1C0BFBEBDBCBBBAB9B8A;
defparam prom_inst_4.INIT_RAM_1D = 256'h827262524232211101F1E1D1C1B1A190807060504030200FFFEFDFCFBFAF9F8F;
defparam prom_inst_4.INIT_RAM_1E = 256'h867565554535251505F5E5D4C4B4A494847464544333231303F3E3D3C3B2A292;
defparam prom_inst_4.INIT_RAM_1F = 256'h897968584838281808F8E8D8C8B7A797877767574737271606F6E6D6C6B6A696;
defparam prom_inst_4.INIT_RAM_20 = 256'h8B7B6B5B4B3B2B1B0BFBEBDACABAAA9A8A7A6A5A4A3A2A1909F9E9D9C9B9A999;
defparam prom_inst_4.INIT_RAM_21 = 256'h8E7E6E5E4D3D2D1D0DFDEDDDCDBDAD9D8D7D6C5C4C3C2C1C0CFCECDCCCBCAC9B;
defparam prom_inst_4.INIT_RAM_22 = 256'h90807060503F2F1F0FFFEFDFCFBFAF9F8F7F6F5F4F3F2E1E0EFEEEDECEBEAE9E;
defparam prom_inst_4.INIT_RAM_23 = 256'h91817161514131211101F1E1D1C1B1A191817160504030201000F0E0D0C0B0A0;
defparam prom_inst_4.INIT_RAM_24 = 256'h93837363534232221202F2E2D2C2B2A292827262524232221202F2E2D2C2B2A1;
defparam prom_inst_4.INIT_RAM_25 = 256'h94847363534333231303F3E3D3C3B3A393837363534333231303F3E3D3C3B3A3;
defparam prom_inst_4.INIT_RAM_26 = 256'h94847464544434241404F4E4D4C4B4A494847464544434241404F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_27 = 256'h94847464544434241404F4E4D4C4B4A494847464544434241404F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_28 = 256'h94847464544434241404F4E4D4C4B4A494847464544434241404F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_29 = 256'h93837363534333231303F3E3D3C3B3A393837363534333231304F4E4D4C4B4A4;
defparam prom_inst_4.INIT_RAM_2A = 256'h92827262524232221202F2E2D2C2B2A292827262524233231303F3E3D3C3B3A3;
defparam prom_inst_4.INIT_RAM_2B = 256'h90807060504030201000F0E1D1C1B1A191817161514131211101F1E1D1C1B2A2;
defparam prom_inst_4.INIT_RAM_2C = 256'h8E7E6E5E4E3E2E1E0EFEEEDFCFBFAF9F8F7F6F5F4F3F2F1F0FFFF0E0D0C0B0A0;
defparam prom_inst_4.INIT_RAM_2D = 256'h8B7B6B5B4C3C2C1C0CFCECDCCCBCAC9C8D7D6D5D4D3D2D1D0DFDEDDDCDBEAE9E;
defparam prom_inst_4.INIT_RAM_2E = 256'h887868584839291909F9E9D9C9B9A99A8A7A6A5A4A3A2A1A0AFBEBDBCBBBAB9B;
defparam prom_inst_4.INIT_RAM_2F = 256'h857565554535251505F6E6D6C6B6A696867667574737271707F7E7D8C8B8A898;
defparam prom_inst_4.INIT_RAM_30 = 256'h807161514131211102F2E2D2C2B2A292837363534333231304F4E4D4C4B4A494;
defparam prom_inst_4.INIT_RAM_31 = 256'h7C6C5C4C3C2D1D0DFDEDDDCEBEAE9E8E7E6E5F4F3F2F1F0FFFF0E0D0C0B0A090;
defparam prom_inst_4.INIT_RAM_32 = 256'h7767574737281808F8E8D8C9B9A99989796A5A4A3A2A1A0BFBEBDBCBBBAB9C8C;
defparam prom_inst_4.INIT_RAM_33 = 256'h7161524232221203F3E3D3C3B3A494847464544535251505F5E6D6C6B6A69687;
defparam prom_inst_4.INIT_RAM_34 = 256'h6B5B4C3C2C1C0CFDEDDDCDBDAD9E8E7E6E5E4F3F2F1F0F00F0E0D0C0B0A19181;
defparam prom_inst_4.INIT_RAM_35 = 256'h64554535251606F6E6D6C7B7A797877868584838291909F9EADACABAAA9B8B7B;
defparam prom_inst_4.INIT_RAM_36 = 256'h5D4E3E2E1E0EFFEFDFCFC0B0A090807161514132221202F2E3D3C3B3A4948474;
defparam prom_inst_4.INIT_RAM_37 = 256'h564636261707F7E7D8C8B8A898897969594A3A2A1A0BFBEBDBCCBCAC9C8D7D6D;
defparam prom_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000E3D3C4B4A495857565;
defparam prom_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[23:0],dout[47:40]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 8;
defparam prom_inst_5.RESET_MODE = "ASYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0C0C0C0C0C;
defparam prom_inst_5.INIT_RAM_01 = 256'h1010101010101010101010100F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0E0E0E0E;
defparam prom_inst_5.INIT_RAM_02 = 256'h1212121212121212121212121211111111111111111111111111111110101010;
defparam prom_inst_5.INIT_RAM_03 = 256'h1414141414141414141414141413131313131313131313131313131313121212;
defparam prom_inst_5.INIT_RAM_04 = 256'h1616161616161616161616161616151515151515151515151515151515151414;
defparam prom_inst_5.INIT_RAM_05 = 256'h1818181818181818181818181818171717171717171717171717171717171616;
defparam prom_inst_5.INIT_RAM_06 = 256'h1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1919191919191919191919191919191918;
defparam prom_inst_5.INIT_RAM_07 = 256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1A;
defparam prom_inst_5.INIT_RAM_08 = 256'h1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D;
defparam prom_inst_5.INIT_RAM_09 = 256'h21202020202020202020202020202020201F1F1F1F1F1F1F1F1F1F1F1F1F1F1F;
defparam prom_inst_5.INIT_RAM_0A = 256'h2322222222222222222222222222222222212121212121212121212121212121;
defparam prom_inst_5.INIT_RAM_0B = 256'h2525242424242424242424242424242424242323232323232323232323232323;
defparam prom_inst_5.INIT_RAM_0C = 256'h2727262626262626262626262626262626262525252525252525252525252525;
defparam prom_inst_5.INIT_RAM_0D = 256'h2929292828282828282828282828282828282827272727272727272727272727;
defparam prom_inst_5.INIT_RAM_0E = 256'h2B2B2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A29292929292929292929292929;
defparam prom_inst_5.INIT_RAM_0F = 256'h2D2D2D2D2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2B2B2B2B2B;
defparam prom_inst_5.INIT_RAM_10 = 256'h2F2F2F2F2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2D2D2D2D2D2D2D2D2D2D2D2D;
defparam prom_inst_5.INIT_RAM_11 = 256'h31313131313030303030303030303030303030302F2F2F2F2F2F2F2F2F2F2F2F;
defparam prom_inst_5.INIT_RAM_12 = 256'h3333333333323232323232323232323232323232323131313131313131313131;
defparam prom_inst_5.INIT_RAM_13 = 256'h3535353535343434343434343434343434343434343333333333333333333333;
defparam prom_inst_5.INIT_RAM_14 = 256'h3737373737373636363636363636363636363636363635353535353535353535;
defparam prom_inst_5.INIT_RAM_15 = 256'h3939393939393838383838383838383838383838383837373737373737373737;
defparam prom_inst_5.INIT_RAM_16 = 256'h3B3B3B3B3B3B3B3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A39393939393939393939;
defparam prom_inst_5.INIT_RAM_17 = 256'h3D3D3D3D3D3D3D3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3B3B3B3B3B3B3B3B3B;
defparam prom_inst_5.INIT_RAM_18 = 256'h3F3F3F3F3F3F3F3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3D3D3D3D3D3D3D3D3D;
defparam prom_inst_5.INIT_RAM_19 = 256'h41414141414141414040404040404040404040404040403F3F3F3F3F3F3F3F3F;
defparam prom_inst_5.INIT_RAM_1A = 256'h4343434343434343424242424242424242424242424242424141414141414141;
defparam prom_inst_5.INIT_RAM_1B = 256'h4545454545454545444444444444444444444444444444444343434343434343;
defparam prom_inst_5.INIT_RAM_1C = 256'h4747474747474747464646464646464646464646464646464545454545454545;
defparam prom_inst_5.INIT_RAM_1D = 256'h4949494949494949494848484848484848484848484848484747474747474747;
defparam prom_inst_5.INIT_RAM_1E = 256'h4B4B4B4B4B4B4B4B4B4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A49494949494949;
defparam prom_inst_5.INIT_RAM_1F = 256'h4D4D4D4D4D4D4D4D4D4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4B4B4B4B4B4B4B;
defparam prom_inst_5.INIT_RAM_20 = 256'h4F4F4F4F4F4F4F4F4F4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4D4D4D4D4D4D4D;
defparam prom_inst_5.INIT_RAM_21 = 256'h515151515151515151505050505050505050505050505050504F4F4F4F4F4F4F;
defparam prom_inst_5.INIT_RAM_22 = 256'h5353535353535353535252525252525252525252525252525251515151515151;
defparam prom_inst_5.INIT_RAM_23 = 256'h5555555555555555555554545454545454545454545454545454535353535353;
defparam prom_inst_5.INIT_RAM_24 = 256'h5757575757575757575756565656565656565656565656565656555555555555;
defparam prom_inst_5.INIT_RAM_25 = 256'h5959595959595959595958585858585858585858585858585858575757575757;
defparam prom_inst_5.INIT_RAM_26 = 256'h5B5B5B5B5B5B5B5B5B5B5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A595959595959;
defparam prom_inst_5.INIT_RAM_27 = 256'h5D5D5D5D5D5D5D5D5D5D5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5B5B5B5B5B5B;
defparam prom_inst_5.INIT_RAM_28 = 256'h5F5F5F5F5F5F5F5F5F5F5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5D5D5D5D5D5D;
defparam prom_inst_5.INIT_RAM_29 = 256'h61616161616161616161606060606060606060606060606060605F5F5F5F5F5F;
defparam prom_inst_5.INIT_RAM_2A = 256'h6363636363636363636362626262626262626262626262626262616161616161;
defparam prom_inst_5.INIT_RAM_2B = 256'h6565656565656565656564646464646464646464646464646464636363636363;
defparam prom_inst_5.INIT_RAM_2C = 256'h6767676767676767676666666666666666666666666666666665656565656565;
defparam prom_inst_5.INIT_RAM_2D = 256'h6969696969696969696868686868686868686868686868686867676767676767;
defparam prom_inst_5.INIT_RAM_2E = 256'h6B6B6B6B6B6B6B6B6B6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A69696969696969;
defparam prom_inst_5.INIT_RAM_2F = 256'h6D6D6D6D6D6D6D6D6D6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6B6B6B6B6B6B6B;
defparam prom_inst_5.INIT_RAM_30 = 256'h6F6F6F6F6F6F6F6F6F6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6D6D6D6D6D6D6D;
defparam prom_inst_5.INIT_RAM_31 = 256'h7171717171717171707070707070707070707070707070706F6F6F6F6F6F6F6F;
defparam prom_inst_5.INIT_RAM_32 = 256'h7373737373737373727272727272727272727272727272727171717171717171;
defparam prom_inst_5.INIT_RAM_33 = 256'h7575757575757575747474747474747474747474747474747373737373737373;
defparam prom_inst_5.INIT_RAM_34 = 256'h7777777777777776767676767676767676767676767676767575757575757575;
defparam prom_inst_5.INIT_RAM_35 = 256'h7979797979797978787878787878787878787878787878777777777777777777;
defparam prom_inst_5.INIT_RAM_36 = 256'h7B7B7B7B7B7B7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A7A797979797979797979;
defparam prom_inst_5.INIT_RAM_37 = 256'h7D7D7D7D7D7D7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7B7B7B7B7B7B7B7B7B7B;
defparam prom_inst_5.INIT_RAM_38 = 256'h00000000000000000000000000000000000000000000007D7D7D7D7D7D7D7D7D;
defparam prom_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //romcoef_module
